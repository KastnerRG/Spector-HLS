
//------> /usr/local/bin/Mentor_Graphics/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /usr/local/bin/Mentor_Graphics/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /usr/local/bin/Mentor_Graphics/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Block 1R1W Read Before Write RAM with common clock
module BLOCK_1R1W_RBW
#(
parameter data_width = 8,
parameter addr_width = 7,
parameter depth = 128
)(
	radr, wadr, d, we, re, clk, q
);

	input [addr_width-1:0] radr;
	input [addr_width-1:0] wadr;
	input [data_width-1:0] d;
	input we;
	input re;
	input clk;
	output[data_width-1:0] q;

	reg [data_width-1:0] q;

	(* ram_style = "block" *)
	reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block_ram"
	//pragma attribute mem block_ram true
		
	always @(posedge clk) begin
		if (we) begin
			mem[wadr] <= d; // Write port
		end
		if (re) begin
			q <= mem[radr] ; // read port
		end
	end

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   mdk@mdk-FX504
//  Generated date: Sat Jan  4 23:55:00 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_7_100_6_gen
// ------------------------------------------------------------------


module SAD_MATCH_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_7_100_6_gen (
  we, d, wadr, re, q, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d
);
  output we;
  output [7:0] d;
  output [6:0] wadr;
  output re;
  input [7:0] q;
  output [6:0] radr;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input [7:0] d_d;
  input we_d;
  input re_d;
  output [7:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_7_100_5_gen
// ------------------------------------------------------------------


module SAD_MATCH_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_7_100_5_gen (
  we, d, wadr, re, q, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d
);
  output we;
  output [7:0] d;
  output [6:0] wadr;
  output re;
  input [7:0] q;
  output [6:0] radr;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input [7:0] d_d;
  input we_d;
  input re_d;
  output [7:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module SAD_MATCH_core_core_fsm (
  clk, rst, core_wen, fsm_output, loop_3_C_2_tr0, loop_2_C_0_tr0, loop_4_C_2_tr0,
      loop_6_C_1_tr0, loop_5_C_0_tr0, loop_lmm_C_2_tr0, loop_8_C_2_tr0, loop_7_C_0_tr0,
      loop_lmm_C_4_tr0
);
  input clk;
  input rst;
  input core_wen;
  output [19:0] fsm_output;
  reg [19:0] fsm_output;
  input loop_3_C_2_tr0;
  input loop_2_C_0_tr0;
  input loop_4_C_2_tr0;
  input loop_6_C_1_tr0;
  input loop_5_C_0_tr0;
  input loop_lmm_C_2_tr0;
  input loop_8_C_2_tr0;
  input loop_7_C_0_tr0;
  input loop_lmm_C_4_tr0;


  // FSM State Type Declaration for SAD_MATCH_core_core_fsm_1
  parameter
    main_C_0 = 5'd0,
    loop_lmm_C_0 = 5'd1,
    loop_lmm_C_1 = 5'd2,
    loop_3_C_0 = 5'd3,
    loop_3_C_1 = 5'd4,
    loop_3_C_2 = 5'd5,
    loop_2_C_0 = 5'd6,
    loop_4_C_0 = 5'd7,
    loop_4_C_1 = 5'd8,
    loop_4_C_2 = 5'd9,
    loop_6_C_0 = 5'd10,
    loop_6_C_1 = 5'd11,
    loop_5_C_0 = 5'd12,
    loop_lmm_C_2 = 5'd13,
    loop_8_C_0 = 5'd14,
    loop_8_C_1 = 5'd15,
    loop_8_C_2 = 5'd16,
    loop_7_C_0 = 5'd17,
    loop_lmm_C_3 = 5'd18,
    loop_lmm_C_4 = 5'd19;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SAD_MATCH_core_core_fsm_1
    case (state_var)
      loop_lmm_C_0 : begin
        fsm_output = 20'b00000000000000000010;
        state_var_NS = loop_lmm_C_1;
      end
      loop_lmm_C_1 : begin
        fsm_output = 20'b00000000000000000100;
        state_var_NS = loop_3_C_0;
      end
      loop_3_C_0 : begin
        fsm_output = 20'b00000000000000001000;
        state_var_NS = loop_3_C_1;
      end
      loop_3_C_1 : begin
        fsm_output = 20'b00000000000000010000;
        state_var_NS = loop_3_C_2;
      end
      loop_3_C_2 : begin
        fsm_output = 20'b00000000000000100000;
        if ( loop_3_C_2_tr0 ) begin
          state_var_NS = loop_2_C_0;
        end
        else begin
          state_var_NS = loop_3_C_0;
        end
      end
      loop_2_C_0 : begin
        fsm_output = 20'b00000000000001000000;
        if ( loop_2_C_0_tr0 ) begin
          state_var_NS = loop_4_C_0;
        end
        else begin
          state_var_NS = loop_3_C_0;
        end
      end
      loop_4_C_0 : begin
        fsm_output = 20'b00000000000010000000;
        state_var_NS = loop_4_C_1;
      end
      loop_4_C_1 : begin
        fsm_output = 20'b00000000000100000000;
        state_var_NS = loop_4_C_2;
      end
      loop_4_C_2 : begin
        fsm_output = 20'b00000000001000000000;
        if ( loop_4_C_2_tr0 ) begin
          state_var_NS = loop_6_C_0;
        end
        else begin
          state_var_NS = loop_4_C_0;
        end
      end
      loop_6_C_0 : begin
        fsm_output = 20'b00000000010000000000;
        state_var_NS = loop_6_C_1;
      end
      loop_6_C_1 : begin
        fsm_output = 20'b00000000100000000000;
        if ( loop_6_C_1_tr0 ) begin
          state_var_NS = loop_5_C_0;
        end
        else begin
          state_var_NS = loop_6_C_0;
        end
      end
      loop_5_C_0 : begin
        fsm_output = 20'b00000001000000000000;
        if ( loop_5_C_0_tr0 ) begin
          state_var_NS = loop_lmm_C_2;
        end
        else begin
          state_var_NS = loop_6_C_0;
        end
      end
      loop_lmm_C_2 : begin
        fsm_output = 20'b00000010000000000000;
        if ( loop_lmm_C_2_tr0 ) begin
          state_var_NS = loop_lmm_C_3;
        end
        else begin
          state_var_NS = loop_8_C_0;
        end
      end
      loop_8_C_0 : begin
        fsm_output = 20'b00000100000000000000;
        state_var_NS = loop_8_C_1;
      end
      loop_8_C_1 : begin
        fsm_output = 20'b00001000000000000000;
        state_var_NS = loop_8_C_2;
      end
      loop_8_C_2 : begin
        fsm_output = 20'b00010000000000000000;
        if ( loop_8_C_2_tr0 ) begin
          state_var_NS = loop_7_C_0;
        end
        else begin
          state_var_NS = loop_8_C_0;
        end
      end
      loop_7_C_0 : begin
        fsm_output = 20'b00100000000000000000;
        if ( loop_7_C_0_tr0 ) begin
          state_var_NS = loop_lmm_C_3;
        end
        else begin
          state_var_NS = loop_8_C_0;
        end
      end
      loop_lmm_C_3 : begin
        fsm_output = 20'b01000000000000000000;
        state_var_NS = loop_lmm_C_4;
      end
      loop_lmm_C_4 : begin
        fsm_output = 20'b10000000000000000000;
        if ( loop_lmm_C_4_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = loop_lmm_C_0;
        end
      end
      // main_C_0
      default : begin
        fsm_output = 20'b00000000000000000001;
        state_var_NS = loop_lmm_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_staller
// ------------------------------------------------------------------


module SAD_MATCH_core_staller (
  clk, rst, core_wen, core_wten, INPUT_rsci_wen_comp, OUTPUT_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input INPUT_rsci_wen_comp;
  input OUTPUT_rsci_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = INPUT_rsci_wen_comp & OUTPUT_rsci_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_win_buf_rsci_1_win_buf_rsc_wait_dp
// ------------------------------------------------------------------


module SAD_MATCH_core_win_buf_rsci_1_win_buf_rsc_wait_dp (
  clk, rst, win_buf_rsci_radr_d, win_buf_rsci_wadr_d, win_buf_rsci_d_d, win_buf_rsci_q_d,
      win_buf_rsci_radr_d_core, win_buf_rsci_wadr_d_core, win_buf_rsci_d_d_core,
      win_buf_rsci_q_d_mxwt, win_buf_rsci_biwt, win_buf_rsci_bdwt, win_buf_rsci_radr_d_core_sct,
      win_buf_rsci_wadr_d_core_sct_pff
);
  input clk;
  input rst;
  output [6:0] win_buf_rsci_radr_d;
  output [6:0] win_buf_rsci_wadr_d;
  output [7:0] win_buf_rsci_d_d;
  input [7:0] win_buf_rsci_q_d;
  input [6:0] win_buf_rsci_radr_d_core;
  input [6:0] win_buf_rsci_wadr_d_core;
  input [7:0] win_buf_rsci_d_d_core;
  output [7:0] win_buf_rsci_q_d_mxwt;
  input win_buf_rsci_biwt;
  input win_buf_rsci_bdwt;
  input win_buf_rsci_radr_d_core_sct;
  input win_buf_rsci_wadr_d_core_sct_pff;


  // Interconnect Declarations
  reg win_buf_rsci_bcwt;
  reg [7:0] win_buf_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign win_buf_rsci_q_d_mxwt = MUX_v_8_2_2(win_buf_rsci_q_d, win_buf_rsci_q_d_bfwt,
      win_buf_rsci_bcwt);
  assign win_buf_rsci_radr_d = MUX_v_7_2_2(7'b0000000, win_buf_rsci_radr_d_core,
      win_buf_rsci_radr_d_core_sct);
  assign win_buf_rsci_wadr_d = MUX_v_7_2_2(7'b0000000, win_buf_rsci_wadr_d_core,
      win_buf_rsci_wadr_d_core_sct_pff);
  assign win_buf_rsci_d_d = MUX_v_8_2_2(8'b00000000, win_buf_rsci_d_d_core, win_buf_rsci_wadr_d_core_sct_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      win_buf_rsci_bcwt <= 1'b0;
    end
    else begin
      win_buf_rsci_bcwt <= ~((~(win_buf_rsci_bcwt | win_buf_rsci_biwt)) | win_buf_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    win_buf_rsci_q_d_bfwt <= win_buf_rsci_q_d_mxwt;
  end

  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_win_buf_rsci_1_win_buf_rsc_wait_ctrl
// ------------------------------------------------------------------


module SAD_MATCH_core_win_buf_rsci_1_win_buf_rsc_wait_ctrl (
  core_wen, core_wten, win_buf_rsci_oswt, win_buf_rsci_biwt, win_buf_rsci_bdwt, win_buf_rsci_radr_d_core_sct_pff,
      win_buf_rsci_oswt_pff, win_buf_rsci_wadr_d_core_sct_pff, win_buf_rsci_iswt0_1_pff
);
  input core_wen;
  input core_wten;
  input win_buf_rsci_oswt;
  output win_buf_rsci_biwt;
  output win_buf_rsci_bdwt;
  output win_buf_rsci_radr_d_core_sct_pff;
  input win_buf_rsci_oswt_pff;
  output win_buf_rsci_wadr_d_core_sct_pff;
  input win_buf_rsci_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign win_buf_rsci_bdwt = win_buf_rsci_oswt & core_wen;
  assign win_buf_rsci_biwt = (~ core_wten) & win_buf_rsci_oswt;
  assign win_buf_rsci_radr_d_core_sct_pff = win_buf_rsci_oswt_pff & core_wen;
  assign win_buf_rsci_wadr_d_core_sct_pff = win_buf_rsci_iswt0_1_pff & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_row_buf_rsci_1_row_buf_rsc_wait_dp
// ------------------------------------------------------------------


module SAD_MATCH_core_row_buf_rsci_1_row_buf_rsc_wait_dp (
  clk, rst, row_buf_rsci_radr_d, row_buf_rsci_wadr_d, row_buf_rsci_d_d, row_buf_rsci_q_d,
      row_buf_rsci_radr_d_core, row_buf_rsci_wadr_d_core, row_buf_rsci_d_d_core,
      row_buf_rsci_q_d_mxwt, row_buf_rsci_biwt, row_buf_rsci_bdwt, row_buf_rsci_radr_d_core_sct,
      row_buf_rsci_wadr_d_core_sct_pff
);
  input clk;
  input rst;
  output [6:0] row_buf_rsci_radr_d;
  output [6:0] row_buf_rsci_wadr_d;
  output [7:0] row_buf_rsci_d_d;
  input [7:0] row_buf_rsci_q_d;
  input [6:0] row_buf_rsci_radr_d_core;
  input [6:0] row_buf_rsci_wadr_d_core;
  input [7:0] row_buf_rsci_d_d_core;
  output [7:0] row_buf_rsci_q_d_mxwt;
  input row_buf_rsci_biwt;
  input row_buf_rsci_bdwt;
  input row_buf_rsci_radr_d_core_sct;
  input row_buf_rsci_wadr_d_core_sct_pff;


  // Interconnect Declarations
  reg row_buf_rsci_bcwt;
  reg [7:0] row_buf_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign row_buf_rsci_q_d_mxwt = MUX_v_8_2_2(row_buf_rsci_q_d, row_buf_rsci_q_d_bfwt,
      row_buf_rsci_bcwt);
  assign row_buf_rsci_radr_d = MUX_v_7_2_2(7'b0000000, row_buf_rsci_radr_d_core,
      row_buf_rsci_radr_d_core_sct);
  assign row_buf_rsci_wadr_d = MUX_v_7_2_2(7'b0000000, row_buf_rsci_wadr_d_core,
      row_buf_rsci_wadr_d_core_sct_pff);
  assign row_buf_rsci_d_d = MUX_v_8_2_2(8'b00000000, row_buf_rsci_d_d_core, row_buf_rsci_wadr_d_core_sct_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      row_buf_rsci_bcwt <= 1'b0;
    end
    else begin
      row_buf_rsci_bcwt <= ~((~(row_buf_rsci_bcwt | row_buf_rsci_biwt)) | row_buf_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    row_buf_rsci_q_d_bfwt <= row_buf_rsci_q_d_mxwt;
  end

  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_row_buf_rsci_1_row_buf_rsc_wait_ctrl
// ------------------------------------------------------------------


module SAD_MATCH_core_row_buf_rsci_1_row_buf_rsc_wait_ctrl (
  core_wen, core_wten, row_buf_rsci_oswt, row_buf_rsci_biwt, row_buf_rsci_bdwt, row_buf_rsci_radr_d_core_sct_pff,
      row_buf_rsci_oswt_pff, row_buf_rsci_wadr_d_core_sct_pff, row_buf_rsci_iswt0_1_pff
);
  input core_wen;
  input core_wten;
  input row_buf_rsci_oswt;
  output row_buf_rsci_biwt;
  output row_buf_rsci_bdwt;
  output row_buf_rsci_radr_d_core_sct_pff;
  input row_buf_rsci_oswt_pff;
  output row_buf_rsci_wadr_d_core_sct_pff;
  input row_buf_rsci_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign row_buf_rsci_bdwt = row_buf_rsci_oswt & core_wen;
  assign row_buf_rsci_biwt = (~ core_wten) & row_buf_rsci_oswt;
  assign row_buf_rsci_radr_d_core_sct_pff = row_buf_rsci_oswt_pff & core_wen;
  assign row_buf_rsci_wadr_d_core_sct_pff = row_buf_rsci_iswt0_1_pff & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_OUTPUT_rsci_OUTPUT_wait_dp
// ------------------------------------------------------------------


module SAD_MATCH_core_OUTPUT_rsci_OUTPUT_wait_dp (
  clk, rst, OUTPUT_rsci_oswt, OUTPUT_rsci_wen_comp, OUTPUT_rsci_biwt, OUTPUT_rsci_bdwt,
      OUTPUT_rsci_bcwt
);
  input clk;
  input rst;
  input OUTPUT_rsci_oswt;
  output OUTPUT_rsci_wen_comp;
  input OUTPUT_rsci_biwt;
  input OUTPUT_rsci_bdwt;
  output OUTPUT_rsci_bcwt;
  reg OUTPUT_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign OUTPUT_rsci_wen_comp = (~ OUTPUT_rsci_oswt) | OUTPUT_rsci_biwt | OUTPUT_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      OUTPUT_rsci_bcwt <= 1'b0;
    end
    else begin
      OUTPUT_rsci_bcwt <= ~((~(OUTPUT_rsci_bcwt | OUTPUT_rsci_biwt)) | OUTPUT_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_OUTPUT_rsci_OUTPUT_wait_ctrl
// ------------------------------------------------------------------


module SAD_MATCH_core_OUTPUT_rsci_OUTPUT_wait_ctrl (
  core_wen, OUTPUT_rsci_oswt, OUTPUT_rsci_irdy, OUTPUT_rsci_biwt, OUTPUT_rsci_bdwt,
      OUTPUT_rsci_bcwt, OUTPUT_rsci_ivld_core_sct
);
  input core_wen;
  input OUTPUT_rsci_oswt;
  input OUTPUT_rsci_irdy;
  output OUTPUT_rsci_biwt;
  output OUTPUT_rsci_bdwt;
  input OUTPUT_rsci_bcwt;
  output OUTPUT_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire OUTPUT_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign OUTPUT_rsci_bdwt = OUTPUT_rsci_oswt & core_wen;
  assign OUTPUT_rsci_biwt = OUTPUT_rsci_ogwt & OUTPUT_rsci_irdy;
  assign OUTPUT_rsci_ogwt = OUTPUT_rsci_oswt & (~ OUTPUT_rsci_bcwt);
  assign OUTPUT_rsci_ivld_core_sct = OUTPUT_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_INPUT_rsci_INPUT_wait_dp
// ------------------------------------------------------------------


module SAD_MATCH_core_INPUT_rsci_INPUT_wait_dp (
  clk, rst, INPUT_rsci_oswt, INPUT_rsci_wen_comp, INPUT_rsci_idat_mxwt, INPUT_rsci_biwt,
      INPUT_rsci_bdwt, INPUT_rsci_bcwt, INPUT_rsci_idat
);
  input clk;
  input rst;
  input INPUT_rsci_oswt;
  output INPUT_rsci_wen_comp;
  output [7:0] INPUT_rsci_idat_mxwt;
  input INPUT_rsci_biwt;
  input INPUT_rsci_bdwt;
  output INPUT_rsci_bcwt;
  reg INPUT_rsci_bcwt;
  input [7:0] INPUT_rsci_idat;


  // Interconnect Declarations
  reg [7:0] INPUT_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign INPUT_rsci_wen_comp = (~ INPUT_rsci_oswt) | INPUT_rsci_biwt | INPUT_rsci_bcwt;
  assign INPUT_rsci_idat_mxwt = MUX_v_8_2_2(INPUT_rsci_idat, INPUT_rsci_idat_bfwt,
      INPUT_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      INPUT_rsci_bcwt <= 1'b0;
    end
    else begin
      INPUT_rsci_bcwt <= ~((~(INPUT_rsci_bcwt | INPUT_rsci_biwt)) | INPUT_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    INPUT_rsci_idat_bfwt <= INPUT_rsci_idat_mxwt;
  end

  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_INPUT_rsci_INPUT_wait_ctrl
// ------------------------------------------------------------------


module SAD_MATCH_core_INPUT_rsci_INPUT_wait_ctrl (
  core_wen, INPUT_rsci_oswt, INPUT_rsci_biwt, INPUT_rsci_bdwt, INPUT_rsci_bcwt, INPUT_rsci_irdy_core_sct,
      INPUT_rsci_ivld
);
  input core_wen;
  input INPUT_rsci_oswt;
  output INPUT_rsci_biwt;
  output INPUT_rsci_bdwt;
  input INPUT_rsci_bcwt;
  output INPUT_rsci_irdy_core_sct;
  input INPUT_rsci_ivld;


  // Interconnect Declarations
  wire INPUT_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign INPUT_rsci_bdwt = INPUT_rsci_oswt & core_wen;
  assign INPUT_rsci_biwt = INPUT_rsci_ogwt & INPUT_rsci_ivld;
  assign INPUT_rsci_ogwt = INPUT_rsci_oswt & (~ INPUT_rsci_bcwt);
  assign INPUT_rsci_irdy_core_sct = INPUT_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_win_buf_rsci_1
// ------------------------------------------------------------------


module SAD_MATCH_core_win_buf_rsci_1 (
  clk, rst, win_buf_rsci_radr_d, win_buf_rsci_wadr_d, win_buf_rsci_d_d, win_buf_rsci_we_d,
      win_buf_rsci_re_d, win_buf_rsci_q_d, core_wen, core_wten, win_buf_rsci_oswt,
      win_buf_rsci_radr_d_core, win_buf_rsci_wadr_d_core, win_buf_rsci_d_d_core,
      win_buf_rsci_q_d_mxwt, win_buf_rsci_oswt_pff, win_buf_rsci_iswt0_1_pff
);
  input clk;
  input rst;
  output [6:0] win_buf_rsci_radr_d;
  output [6:0] win_buf_rsci_wadr_d;
  output [7:0] win_buf_rsci_d_d;
  output win_buf_rsci_we_d;
  output win_buf_rsci_re_d;
  input [7:0] win_buf_rsci_q_d;
  input core_wen;
  input core_wten;
  input win_buf_rsci_oswt;
  input [6:0] win_buf_rsci_radr_d_core;
  input [6:0] win_buf_rsci_wadr_d_core;
  input [7:0] win_buf_rsci_d_d_core;
  output [7:0] win_buf_rsci_q_d_mxwt;
  input win_buf_rsci_oswt_pff;
  input win_buf_rsci_iswt0_1_pff;


  // Interconnect Declarations
  wire win_buf_rsci_biwt;
  wire win_buf_rsci_bdwt;
  wire [6:0] win_buf_rsci_radr_d_reg;
  wire win_buf_rsci_radr_d_core_sct_iff;
  wire [6:0] win_buf_rsci_wadr_d_reg;
  wire win_buf_rsci_wadr_d_core_sct_iff;
  wire [7:0] win_buf_rsci_d_d_reg;


  // Interconnect Declarations for Component Instantiations 
  SAD_MATCH_core_win_buf_rsci_1_win_buf_rsc_wait_ctrl SAD_MATCH_core_win_buf_rsci_1_win_buf_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .win_buf_rsci_oswt(win_buf_rsci_oswt),
      .win_buf_rsci_biwt(win_buf_rsci_biwt),
      .win_buf_rsci_bdwt(win_buf_rsci_bdwt),
      .win_buf_rsci_radr_d_core_sct_pff(win_buf_rsci_radr_d_core_sct_iff),
      .win_buf_rsci_oswt_pff(win_buf_rsci_oswt_pff),
      .win_buf_rsci_wadr_d_core_sct_pff(win_buf_rsci_wadr_d_core_sct_iff),
      .win_buf_rsci_iswt0_1_pff(win_buf_rsci_iswt0_1_pff)
    );
  SAD_MATCH_core_win_buf_rsci_1_win_buf_rsc_wait_dp SAD_MATCH_core_win_buf_rsci_1_win_buf_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .win_buf_rsci_radr_d(win_buf_rsci_radr_d_reg),
      .win_buf_rsci_wadr_d(win_buf_rsci_wadr_d_reg),
      .win_buf_rsci_d_d(win_buf_rsci_d_d_reg),
      .win_buf_rsci_q_d(win_buf_rsci_q_d),
      .win_buf_rsci_radr_d_core(win_buf_rsci_radr_d_core),
      .win_buf_rsci_wadr_d_core(win_buf_rsci_wadr_d_core),
      .win_buf_rsci_d_d_core(win_buf_rsci_d_d_core),
      .win_buf_rsci_q_d_mxwt(win_buf_rsci_q_d_mxwt),
      .win_buf_rsci_biwt(win_buf_rsci_biwt),
      .win_buf_rsci_bdwt(win_buf_rsci_bdwt),
      .win_buf_rsci_radr_d_core_sct(win_buf_rsci_radr_d_core_sct_iff),
      .win_buf_rsci_wadr_d_core_sct_pff(win_buf_rsci_wadr_d_core_sct_iff)
    );
  assign win_buf_rsci_radr_d = win_buf_rsci_radr_d_reg;
  assign win_buf_rsci_wadr_d = win_buf_rsci_wadr_d_reg;
  assign win_buf_rsci_d_d = win_buf_rsci_d_d_reg;
  assign win_buf_rsci_we_d = win_buf_rsci_wadr_d_core_sct_iff;
  assign win_buf_rsci_re_d = win_buf_rsci_radr_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_row_buf_rsci_1
// ------------------------------------------------------------------


module SAD_MATCH_core_row_buf_rsci_1 (
  clk, rst, row_buf_rsci_radr_d, row_buf_rsci_wadr_d, row_buf_rsci_d_d, row_buf_rsci_we_d,
      row_buf_rsci_re_d, row_buf_rsci_q_d, core_wen, core_wten, row_buf_rsci_oswt,
      row_buf_rsci_radr_d_core, row_buf_rsci_wadr_d_core, row_buf_rsci_d_d_core,
      row_buf_rsci_q_d_mxwt, row_buf_rsci_oswt_pff, row_buf_rsci_iswt0_1_pff
);
  input clk;
  input rst;
  output [6:0] row_buf_rsci_radr_d;
  output [6:0] row_buf_rsci_wadr_d;
  output [7:0] row_buf_rsci_d_d;
  output row_buf_rsci_we_d;
  output row_buf_rsci_re_d;
  input [7:0] row_buf_rsci_q_d;
  input core_wen;
  input core_wten;
  input row_buf_rsci_oswt;
  input [6:0] row_buf_rsci_radr_d_core;
  input [6:0] row_buf_rsci_wadr_d_core;
  input [7:0] row_buf_rsci_d_d_core;
  output [7:0] row_buf_rsci_q_d_mxwt;
  input row_buf_rsci_oswt_pff;
  input row_buf_rsci_iswt0_1_pff;


  // Interconnect Declarations
  wire row_buf_rsci_biwt;
  wire row_buf_rsci_bdwt;
  wire [6:0] row_buf_rsci_radr_d_reg;
  wire row_buf_rsci_radr_d_core_sct_iff;
  wire [6:0] row_buf_rsci_wadr_d_reg;
  wire row_buf_rsci_wadr_d_core_sct_iff;
  wire [7:0] row_buf_rsci_d_d_reg;


  // Interconnect Declarations for Component Instantiations 
  SAD_MATCH_core_row_buf_rsci_1_row_buf_rsc_wait_ctrl SAD_MATCH_core_row_buf_rsci_1_row_buf_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .row_buf_rsci_oswt(row_buf_rsci_oswt),
      .row_buf_rsci_biwt(row_buf_rsci_biwt),
      .row_buf_rsci_bdwt(row_buf_rsci_bdwt),
      .row_buf_rsci_radr_d_core_sct_pff(row_buf_rsci_radr_d_core_sct_iff),
      .row_buf_rsci_oswt_pff(row_buf_rsci_oswt_pff),
      .row_buf_rsci_wadr_d_core_sct_pff(row_buf_rsci_wadr_d_core_sct_iff),
      .row_buf_rsci_iswt0_1_pff(row_buf_rsci_iswt0_1_pff)
    );
  SAD_MATCH_core_row_buf_rsci_1_row_buf_rsc_wait_dp SAD_MATCH_core_row_buf_rsci_1_row_buf_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .row_buf_rsci_radr_d(row_buf_rsci_radr_d_reg),
      .row_buf_rsci_wadr_d(row_buf_rsci_wadr_d_reg),
      .row_buf_rsci_d_d(row_buf_rsci_d_d_reg),
      .row_buf_rsci_q_d(row_buf_rsci_q_d),
      .row_buf_rsci_radr_d_core(row_buf_rsci_radr_d_core),
      .row_buf_rsci_wadr_d_core(row_buf_rsci_wadr_d_core),
      .row_buf_rsci_d_d_core(row_buf_rsci_d_d_core),
      .row_buf_rsci_q_d_mxwt(row_buf_rsci_q_d_mxwt),
      .row_buf_rsci_biwt(row_buf_rsci_biwt),
      .row_buf_rsci_bdwt(row_buf_rsci_bdwt),
      .row_buf_rsci_radr_d_core_sct(row_buf_rsci_radr_d_core_sct_iff),
      .row_buf_rsci_wadr_d_core_sct_pff(row_buf_rsci_wadr_d_core_sct_iff)
    );
  assign row_buf_rsci_radr_d = row_buf_rsci_radr_d_reg;
  assign row_buf_rsci_wadr_d = row_buf_rsci_wadr_d_reg;
  assign row_buf_rsci_d_d = row_buf_rsci_d_d_reg;
  assign row_buf_rsci_we_d = row_buf_rsci_wadr_d_core_sct_iff;
  assign row_buf_rsci_re_d = row_buf_rsci_radr_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_OUTPUT_rsci
// ------------------------------------------------------------------


module SAD_MATCH_core_OUTPUT_rsci (
  clk, rst, OUTPUT_rsc_dat, OUTPUT_rsc_vld, OUTPUT_rsc_rdy, core_wen, OUTPUT_rsci_oswt,
      OUTPUT_rsci_wen_comp, OUTPUT_rsci_idat
);
  input clk;
  input rst;
  output [7:0] OUTPUT_rsc_dat;
  output OUTPUT_rsc_vld;
  input OUTPUT_rsc_rdy;
  input core_wen;
  input OUTPUT_rsci_oswt;
  output OUTPUT_rsci_wen_comp;
  input [7:0] OUTPUT_rsci_idat;


  // Interconnect Declarations
  wire OUTPUT_rsci_irdy;
  wire OUTPUT_rsci_biwt;
  wire OUTPUT_rsci_bdwt;
  wire OUTPUT_rsci_bcwt;
  wire OUTPUT_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_OUTPUT_rsci_idat;
  assign nl_OUTPUT_rsci_idat = {7'b0000000 , (OUTPUT_rsci_idat[0])};
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd8)) OUTPUT_rsci (
      .irdy(OUTPUT_rsci_irdy),
      .ivld(OUTPUT_rsci_ivld_core_sct),
      .idat(nl_OUTPUT_rsci_idat[7:0]),
      .rdy(OUTPUT_rsc_rdy),
      .vld(OUTPUT_rsc_vld),
      .dat(OUTPUT_rsc_dat)
    );
  SAD_MATCH_core_OUTPUT_rsci_OUTPUT_wait_ctrl SAD_MATCH_core_OUTPUT_rsci_OUTPUT_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .OUTPUT_rsci_oswt(OUTPUT_rsci_oswt),
      .OUTPUT_rsci_irdy(OUTPUT_rsci_irdy),
      .OUTPUT_rsci_biwt(OUTPUT_rsci_biwt),
      .OUTPUT_rsci_bdwt(OUTPUT_rsci_bdwt),
      .OUTPUT_rsci_bcwt(OUTPUT_rsci_bcwt),
      .OUTPUT_rsci_ivld_core_sct(OUTPUT_rsci_ivld_core_sct)
    );
  SAD_MATCH_core_OUTPUT_rsci_OUTPUT_wait_dp SAD_MATCH_core_OUTPUT_rsci_OUTPUT_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .OUTPUT_rsci_oswt(OUTPUT_rsci_oswt),
      .OUTPUT_rsci_wen_comp(OUTPUT_rsci_wen_comp),
      .OUTPUT_rsci_biwt(OUTPUT_rsci_biwt),
      .OUTPUT_rsci_bdwt(OUTPUT_rsci_bdwt),
      .OUTPUT_rsci_bcwt(OUTPUT_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core_INPUT_rsci
// ------------------------------------------------------------------


module SAD_MATCH_core_INPUT_rsci (
  clk, rst, INPUT_rsc_dat, INPUT_rsc_vld, INPUT_rsc_rdy, core_wen, INPUT_rsci_oswt,
      INPUT_rsci_wen_comp, INPUT_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [7:0] INPUT_rsc_dat;
  input INPUT_rsc_vld;
  output INPUT_rsc_rdy;
  input core_wen;
  input INPUT_rsci_oswt;
  output INPUT_rsci_wen_comp;
  output [7:0] INPUT_rsci_idat_mxwt;


  // Interconnect Declarations
  wire INPUT_rsci_biwt;
  wire INPUT_rsci_bdwt;
  wire INPUT_rsci_bcwt;
  wire INPUT_rsci_irdy_core_sct;
  wire INPUT_rsci_ivld;
  wire [7:0] INPUT_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd8)) INPUT_rsci (
      .rdy(INPUT_rsc_rdy),
      .vld(INPUT_rsc_vld),
      .dat(INPUT_rsc_dat),
      .irdy(INPUT_rsci_irdy_core_sct),
      .ivld(INPUT_rsci_ivld),
      .idat(INPUT_rsci_idat)
    );
  SAD_MATCH_core_INPUT_rsci_INPUT_wait_ctrl SAD_MATCH_core_INPUT_rsci_INPUT_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .INPUT_rsci_oswt(INPUT_rsci_oswt),
      .INPUT_rsci_biwt(INPUT_rsci_biwt),
      .INPUT_rsci_bdwt(INPUT_rsci_bdwt),
      .INPUT_rsci_bcwt(INPUT_rsci_bcwt),
      .INPUT_rsci_irdy_core_sct(INPUT_rsci_irdy_core_sct),
      .INPUT_rsci_ivld(INPUT_rsci_ivld)
    );
  SAD_MATCH_core_INPUT_rsci_INPUT_wait_dp SAD_MATCH_core_INPUT_rsci_INPUT_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .INPUT_rsci_oswt(INPUT_rsci_oswt),
      .INPUT_rsci_wen_comp(INPUT_rsci_wen_comp),
      .INPUT_rsci_idat_mxwt(INPUT_rsci_idat_mxwt),
      .INPUT_rsci_biwt(INPUT_rsci_biwt),
      .INPUT_rsci_bdwt(INPUT_rsci_bdwt),
      .INPUT_rsci_bcwt(INPUT_rsci_bcwt),
      .INPUT_rsci_idat(INPUT_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH_core
// ------------------------------------------------------------------


module SAD_MATCH_core (
  clk, rst, INPUT_rsc_dat, INPUT_rsc_vld, INPUT_rsc_rdy, OUTPUT_rsc_dat, OUTPUT_rsc_vld,
      OUTPUT_rsc_rdy, row_buf_rsci_radr_d, row_buf_rsci_wadr_d, row_buf_rsci_d_d,
      row_buf_rsci_we_d, row_buf_rsci_re_d, row_buf_rsci_q_d, win_buf_rsci_radr_d,
      win_buf_rsci_wadr_d, win_buf_rsci_d_d, win_buf_rsci_we_d, win_buf_rsci_re_d,
      win_buf_rsci_q_d
);
  input clk;
  input rst;
  input [7:0] INPUT_rsc_dat;
  input INPUT_rsc_vld;
  output INPUT_rsc_rdy;
  output [7:0] OUTPUT_rsc_dat;
  output OUTPUT_rsc_vld;
  input OUTPUT_rsc_rdy;
  output [6:0] row_buf_rsci_radr_d;
  output [6:0] row_buf_rsci_wadr_d;
  output [7:0] row_buf_rsci_d_d;
  output row_buf_rsci_we_d;
  output row_buf_rsci_re_d;
  input [7:0] row_buf_rsci_q_d;
  output [6:0] win_buf_rsci_radr_d;
  output [6:0] win_buf_rsci_wadr_d;
  output [7:0] win_buf_rsci_d_d;
  output win_buf_rsci_we_d;
  output win_buf_rsci_re_d;
  input [7:0] win_buf_rsci_q_d;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire INPUT_rsci_wen_comp;
  wire [7:0] INPUT_rsci_idat_mxwt;
  wire OUTPUT_rsci_wen_comp;
  wire [7:0] row_buf_rsci_q_d_mxwt;
  wire [7:0] win_buf_rsci_q_d_mxwt;
  reg OUTPUT_rsci_idat_0;
  wire [19:0] fsm_output;
  wire and_dcpl_49;
  wire or_dcpl_81;
  wire or_dcpl_83;
  wire or_dcpl_85;
  wire or_tmp_46;
  reg loop_lmm_loop_lmm_nor_itm;
  reg k_sva_3;
  reg loop_3_slc_loop_3_acc_3_itm;
  wire [31:0] k_sva_1_mx1;
  wire k_sva_1_mx2_3;
  reg reg_INPUT_rsci_oswt_cse;
  reg reg_OUTPUT_rsci_oswt_cse;
  reg reg_row_buf_rsci_oswt_cse;
  reg reg_win_buf_rsci_oswt_cse;
  wire [6:0] row_buf_rsci_radr_d_reg;
  wire or_141_rmff;
  wire [6:0] row_buf_rsci_wadr_d_reg;
  wire [7:0] row_buf_rsci_d_d_reg;
  wire row_buf_rsci_we_d_reg;
  wire row_buf_rsci_re_d_reg;
  wire [6:0] win_buf_rsci_radr_d_reg;
  wire [6:0] win_buf_rsci_wadr_d_reg;
  wire [7:0] win_buf_rsci_d_d_reg;
  wire win_buf_rsci_we_d_reg;
  wire win_buf_rsci_re_d_reg;
  reg [3:0] j_3_0_sva;
  reg [1:0] k_sva_7_6;
  reg [1:0] k_sva_5_4;
  reg [5:0] loop_8_acc_10_itm;
  reg [23:0] k_sva_31_8;
  reg [3:0] loop_1_z_3_0_sva;
  reg [3:0] loop_3_acc_14_psp;
  reg [3:0] loop_3_acc_12_sdt_3_0;
  wire [3:0] loop_3_acc_11_sdt_3_0_1;
  wire [4:0] nl_loop_3_acc_11_sdt_3_0_1;
  wire [3:0] z_out;
  wire [4:0] nl_z_out;
  wire or_tmp_86;
  wire [7:0] z_out_3;
  wire [8:0] nl_z_out_3;
  wire or_tmp_89;
  wire [32:0] z_out_4;
  wire [33:0] nl_z_out_4;
  wire [15:0] z_out_6;
  wire [16:0] nl_z_out_6;
  wire [5:0] z_out_7;
  wire [6:0] nl_z_out_7;
  reg [15:0] loop_lmm_i_15_0_sva;
  reg [15:0] i_15_0_sva;
  reg [15:0] loop_op_i_15_0_sva;
  reg [31:0] loop_1_sad_lpi_4;
  reg [31:0] k_sva_1;
  reg [7:0] o_7_0_sva_1;
  wire [15:0] i_15_0_sva_2;
  wire [16:0] nl_i_15_0_sva_2;
  wire j_3_0_sva_mx0c1;
  wire j_3_0_sva_mx0c2;
  wire loop_1_loop_1_nand_seb_1;
  wire loop_1_or_3_ssc;
  wire loop_8_or_ssc;
  wire and_cse;
  wire [15:0] loop_1_loop_1_and_2_cse;
  wire or_218_ssc;
  wire z_out_1_3;
  wire [3:0] z_out_2_3_0;
  wire [31:0] z_out_5_31_0;
  wire [32:0] nl_z_out_5_31_0;

  wire[0:0] loop_op_i_not_nl;
  wire[0:0] not_111_nl;
  wire[23:0] k_mux_5_nl;
  wire[7:0] loop_8_loop_8_and_nl;
  wire[7:0] loop_8_mux_1_nl;
  wire[0:0] or_211_nl;
  wire[0:0] k_not_nl;
  wire[1:0] k_mux_4_nl;
  wire[0:0] nor_29_nl;
  wire[0:0] nor_37_nl;
  wire[0:0] k_mux1h_10_nl;
  wire[0:0] loop_1_loop_1_and_nl;
  wire[0:0] and_146_nl;
  wire[2:0] k_k_and_nl;
  wire[2:0] k_mux_3_nl;
  wire[0:0] nor_32_nl;
  wire[0:0] nor_31_nl;
  wire[3:0] loop_1_z_mux_nl;
  wire[0:0] j_not_nl;
  wire[3:0] n_mux1h_nl;
  wire[0:0] or_163_nl;
  wire[0:0] nor_nl;
  wire[10:0] loop_lmm_acc_nl;
  wire[11:0] nl_loop_lmm_acc_nl;
  wire[10:0] loop_op_acc_nl;
  wire[11:0] nl_loop_op_acc_nl;
  wire[3:0] loop_3_mux_5_nl;
  wire[0:0] loop_3_or_4_nl;
  wire[1:0] loop_3_loop_3_mux_1_nl;
  wire[0:0] loop_3_mux_6_nl;
  wire[0:0] loop_3_mux_7_nl;
  wire[0:0] loop_3_mux_8_nl;
  wire[4:0] acc_2_nl;
  wire[5:0] nl_acc_2_nl;
  wire[3:0] loop_4_mux_1_nl;
  wire[0:0] loop_4_or_1_nl;
  wire[2:0] loop_4_mux1h_1_nl;
  wire[7:0] loop_8_mux_7_nl;
  wire[3:0] loop_8_mux_8_nl;
  wire[31:0] loop_1_mux1h_4_nl;
  wire[0:0] loop_1_or_4_nl;
  wire[0:0] loop_1_or_5_nl;
  wire[8:0] loop_1_or_6_nl;
  wire[0:0] loop_1_loop_1_or_1_nl;
  wire[7:0] loop_1_mux1h_5_nl;
  wire[31:0] loop_8_mux1h_4_nl;
  wire[0:0] loop_8_loop_8_or_3_nl;
  wire[1:0] loop_8_loop_8_or_4_nl;
  wire[0:0] loop_8_not_4_nl;
  wire[1:0] loop_8_loop_8_or_5_nl;
  wire[0:0] loop_8_not_5_nl;
  wire[15:0] loop_lmm_mux_3_nl;
  wire[5:0] loop_8_mux_9_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SAD_MATCH_core_OUTPUT_rsci_inst_OUTPUT_rsci_idat;
  assign nl_SAD_MATCH_core_OUTPUT_rsci_inst_OUTPUT_rsci_idat = {7'b0, OUTPUT_rsci_idat_0};
  wire[5:0] row_buf_mux_1_nl;
  wire[5:0] loop_8_acc_9_nl;
  wire[6:0] nl_loop_8_acc_9_nl;
  wire[5:0] loop_8_acc_12_nl;
  wire[6:0] nl_loop_8_acc_12_nl;
  wire[0:0] row_buf_mux_nl;
  wire [6:0] nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_radr_d_core;
  assign nl_loop_8_acc_12_nl = ({j_3_0_sva , 2'b01}) + conv_u2u_4_6({(z_out_4[1:0])
      , (j_3_0_sva[1:0])});
  assign loop_8_acc_12_nl = nl_loop_8_acc_12_nl[5:0];
  assign nl_loop_8_acc_9_nl = (loop_8_acc_12_nl) + (k_sva_31_8[6:1]);
  assign loop_8_acc_9_nl = nl_loop_8_acc_9_nl[5:0];
  assign row_buf_mux_1_nl = MUX_v_6_2_2(z_out_7, (loop_8_acc_9_nl), fsm_output[14]);
  assign row_buf_mux_nl = MUX_s_1_2_2((loop_8_acc_10_itm[0]), (k_sva_31_8[0]), fsm_output[14]);
  assign nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_radr_d_core = {(row_buf_mux_1_nl)
      , (row_buf_mux_nl)};
  wire[5:0] row_buf_mux_3_nl;
  wire[0:0] row_buf_mux_2_nl;
  wire [6:0] nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_wadr_d_core;
  assign row_buf_mux_3_nl = MUX_v_6_2_2((z_out_4[5:0]), loop_8_acc_10_itm, fsm_output[15]);
  assign row_buf_mux_2_nl = MUX_s_1_2_2((loop_8_acc_10_itm[0]), (k_sva_31_8[0]),
      fsm_output[15]);
  assign nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_wadr_d_core = {(row_buf_mux_3_nl)
      , (row_buf_mux_2_nl)};
  wire [7:0] nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_d_d_core;
  assign nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_d_d_core = MUX_v_8_2_2(INPUT_rsci_idat_mxwt,
      row_buf_rsci_q_d_mxwt, fsm_output[15]);
  wire [0:0] nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_iswt0_1_pff;
  assign nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_iswt0_1_pff = (fsm_output[1])
      | (fsm_output[15]);
  wire[3:0] win_buf_mux_2_nl;
  wire[3:0] loop_3_acc_13_nl;
  wire[4:0] nl_loop_3_acc_13_nl;
  wire[1:0] win_buf_mux_1_nl;
  wire[0:0] win_buf_mux_nl;
  wire [6:0] nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_radr_d_core;
  assign nl_loop_3_acc_13_nl = conv_u2u_2_4(loop_3_acc_11_sdt_3_0_1[3:2]) + loop_1_z_3_0_sva;
  assign loop_3_acc_13_nl = nl_loop_3_acc_13_nl[3:0];
  assign win_buf_mux_2_nl = MUX_v_4_2_2((loop_3_acc_13_nl), z_out, fsm_output[10]);
  assign win_buf_mux_1_nl = MUX_v_2_2_2((loop_3_acc_11_sdt_3_0_1[1:0]), (z_out_2_3_0[1:0]),
      fsm_output[10]);
  assign win_buf_mux_nl = MUX_s_1_2_2((z_out_4[0]), (loop_1_z_3_0_sva[0]), fsm_output[10]);
  assign nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_radr_d_core = {(win_buf_mux_2_nl)
      , (win_buf_mux_1_nl) , (win_buf_mux_nl)};
  wire[3:0] loop_3_mux_nl;
  wire[1:0] win_buf_mux_3_nl;
  wire[0:0] win_buf_win_buf_or_nl;
  wire [6:0] nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_wadr_d_core;
  assign loop_3_mux_nl = MUX_v_4_2_2(loop_3_acc_14_psp, loop_3_acc_12_sdt_3_0, fsm_output[8]);
  assign win_buf_mux_3_nl = MUX_v_2_2_2((loop_3_acc_12_sdt_3_0[1:0]), (j_3_0_sva[1:0]),
      fsm_output[8]);
  assign win_buf_win_buf_or_nl = (j_3_0_sva[0]) | (~ (fsm_output[4]));
  assign nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_wadr_d_core = {(loop_3_mux_nl)
      , (win_buf_mux_3_nl) , (win_buf_win_buf_or_nl)};
  wire [7:0] nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_d_d_core;
  assign nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_d_d_core = MUX_v_8_2_2(win_buf_rsci_q_d_mxwt,
      row_buf_rsci_q_d_mxwt, fsm_output[8]);
  wire [0:0] nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_iswt0_1_pff;
  assign nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_iswt0_1_pff = (fsm_output[8])
      | (fsm_output[4]);
  wire [0:0] nl_SAD_MATCH_core_core_fsm_inst_loop_3_C_2_tr0;
  assign nl_SAD_MATCH_core_core_fsm_inst_loop_3_C_2_tr0 = ~ loop_3_slc_loop_3_acc_3_itm;
  wire [0:0] nl_SAD_MATCH_core_core_fsm_inst_loop_2_C_0_tr0;
  assign nl_SAD_MATCH_core_core_fsm_inst_loop_2_C_0_tr0 = ~ (z_out_3[4]);
  wire [0:0] nl_SAD_MATCH_core_core_fsm_inst_loop_4_C_2_tr0;
  assign nl_SAD_MATCH_core_core_fsm_inst_loop_4_C_2_tr0 = ~ loop_3_slc_loop_3_acc_3_itm;
  wire [0:0] nl_SAD_MATCH_core_core_fsm_inst_loop_6_C_1_tr0;
  assign nl_SAD_MATCH_core_core_fsm_inst_loop_6_C_1_tr0 = ~ loop_3_slc_loop_3_acc_3_itm;
  wire [0:0] nl_SAD_MATCH_core_core_fsm_inst_loop_5_C_0_tr0;
  assign nl_SAD_MATCH_core_core_fsm_inst_loop_5_C_0_tr0 = ~ z_out_1_3;
  wire [0:0] nl_SAD_MATCH_core_core_fsm_inst_loop_lmm_C_2_tr0;
  assign nl_SAD_MATCH_core_core_fsm_inst_loop_lmm_C_2_tr0 = (z_out_5_31_0!=32'b00000000000000000000000011001000);
  wire [0:0] nl_SAD_MATCH_core_core_fsm_inst_loop_8_C_2_tr0;
  assign nl_SAD_MATCH_core_core_fsm_inst_loop_8_C_2_tr0 = ~ k_sva_3;
  wire [0:0] nl_SAD_MATCH_core_core_fsm_inst_loop_7_C_0_tr0;
  assign nl_SAD_MATCH_core_core_fsm_inst_loop_7_C_0_tr0 = ~ (z_out_3[4]);
  SAD_MATCH_core_INPUT_rsci SAD_MATCH_core_INPUT_rsci_inst (
      .clk(clk),
      .rst(rst),
      .INPUT_rsc_dat(INPUT_rsc_dat),
      .INPUT_rsc_vld(INPUT_rsc_vld),
      .INPUT_rsc_rdy(INPUT_rsc_rdy),
      .core_wen(core_wen),
      .INPUT_rsci_oswt(reg_INPUT_rsci_oswt_cse),
      .INPUT_rsci_wen_comp(INPUT_rsci_wen_comp),
      .INPUT_rsci_idat_mxwt(INPUT_rsci_idat_mxwt)
    );
  SAD_MATCH_core_OUTPUT_rsci SAD_MATCH_core_OUTPUT_rsci_inst (
      .clk(clk),
      .rst(rst),
      .OUTPUT_rsc_dat(OUTPUT_rsc_dat),
      .OUTPUT_rsc_vld(OUTPUT_rsc_vld),
      .OUTPUT_rsc_rdy(OUTPUT_rsc_rdy),
      .core_wen(core_wen),
      .OUTPUT_rsci_oswt(reg_OUTPUT_rsci_oswt_cse),
      .OUTPUT_rsci_wen_comp(OUTPUT_rsci_wen_comp),
      .OUTPUT_rsci_idat(nl_SAD_MATCH_core_OUTPUT_rsci_inst_OUTPUT_rsci_idat[7:0])
    );
  SAD_MATCH_core_row_buf_rsci_1 SAD_MATCH_core_row_buf_rsci_1_inst (
      .clk(clk),
      .rst(rst),
      .row_buf_rsci_radr_d(row_buf_rsci_radr_d_reg),
      .row_buf_rsci_wadr_d(row_buf_rsci_wadr_d_reg),
      .row_buf_rsci_d_d(row_buf_rsci_d_d_reg),
      .row_buf_rsci_we_d(row_buf_rsci_we_d_reg),
      .row_buf_rsci_re_d(row_buf_rsci_re_d_reg),
      .row_buf_rsci_q_d(row_buf_rsci_q_d),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .row_buf_rsci_oswt(reg_row_buf_rsci_oswt_cse),
      .row_buf_rsci_radr_d_core(nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_radr_d_core[6:0]),
      .row_buf_rsci_wadr_d_core(nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_wadr_d_core[6:0]),
      .row_buf_rsci_d_d_core(nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_d_d_core[7:0]),
      .row_buf_rsci_q_d_mxwt(row_buf_rsci_q_d_mxwt),
      .row_buf_rsci_oswt_pff(or_141_rmff),
      .row_buf_rsci_iswt0_1_pff(nl_SAD_MATCH_core_row_buf_rsci_1_inst_row_buf_rsci_iswt0_1_pff[0:0])
    );
  SAD_MATCH_core_win_buf_rsci_1 SAD_MATCH_core_win_buf_rsci_1_inst (
      .clk(clk),
      .rst(rst),
      .win_buf_rsci_radr_d(win_buf_rsci_radr_d_reg),
      .win_buf_rsci_wadr_d(win_buf_rsci_wadr_d_reg),
      .win_buf_rsci_d_d(win_buf_rsci_d_d_reg),
      .win_buf_rsci_we_d(win_buf_rsci_we_d_reg),
      .win_buf_rsci_re_d(win_buf_rsci_re_d_reg),
      .win_buf_rsci_q_d(win_buf_rsci_q_d),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .win_buf_rsci_oswt(reg_win_buf_rsci_oswt_cse),
      .win_buf_rsci_radr_d_core(nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_radr_d_core[6:0]),
      .win_buf_rsci_wadr_d_core(nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_wadr_d_core[6:0]),
      .win_buf_rsci_d_d_core(nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_d_d_core[7:0]),
      .win_buf_rsci_q_d_mxwt(win_buf_rsci_q_d_mxwt),
      .win_buf_rsci_oswt_pff(or_tmp_46),
      .win_buf_rsci_iswt0_1_pff(nl_SAD_MATCH_core_win_buf_rsci_1_inst_win_buf_rsci_iswt0_1_pff[0:0])
    );
  SAD_MATCH_core_staller SAD_MATCH_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .INPUT_rsci_wen_comp(INPUT_rsci_wen_comp),
      .OUTPUT_rsci_wen_comp(OUTPUT_rsci_wen_comp)
    );
  SAD_MATCH_core_core_fsm SAD_MATCH_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output),
      .loop_3_C_2_tr0(nl_SAD_MATCH_core_core_fsm_inst_loop_3_C_2_tr0[0:0]),
      .loop_2_C_0_tr0(nl_SAD_MATCH_core_core_fsm_inst_loop_2_C_0_tr0[0:0]),
      .loop_4_C_2_tr0(nl_SAD_MATCH_core_core_fsm_inst_loop_4_C_2_tr0[0:0]),
      .loop_6_C_1_tr0(nl_SAD_MATCH_core_core_fsm_inst_loop_6_C_1_tr0[0:0]),
      .loop_5_C_0_tr0(nl_SAD_MATCH_core_core_fsm_inst_loop_5_C_0_tr0[0:0]),
      .loop_lmm_C_2_tr0(nl_SAD_MATCH_core_core_fsm_inst_loop_lmm_C_2_tr0[0:0]),
      .loop_8_C_2_tr0(nl_SAD_MATCH_core_core_fsm_inst_loop_8_C_2_tr0[0:0]),
      .loop_7_C_0_tr0(nl_SAD_MATCH_core_core_fsm_inst_loop_7_C_0_tr0[0:0]),
      .loop_lmm_C_4_tr0(loop_lmm_loop_lmm_nor_itm)
    );
  assign and_cse = ((fsm_output[18]) | (fsm_output[0])) & core_wen;
  assign loop_op_i_not_nl = ~ (fsm_output[0]);
  assign loop_1_loop_1_and_2_cse = MUX_v_16_2_2(16'b0000000000000000, z_out_6, (loop_op_i_not_nl));
  assign or_141_rmff = (fsm_output[7]) | (fsm_output[14]);
  assign nl_i_15_0_sva_2 = i_15_0_sva + 16'b0000000000000001;
  assign i_15_0_sva_2 = nl_i_15_0_sva_2[15:0];
  assign nl_loop_3_acc_11_sdt_3_0_1 = loop_1_z_3_0_sva + conv_u2u_3_4(z_out_4[3:1]);
  assign loop_3_acc_11_sdt_3_0_1 = nl_loop_3_acc_11_sdt_3_0_1[3:0];
  assign k_sva_1_mx1 = MUX_v_32_2_2(k_sva_1, z_out_5_31_0, fsm_output[13]);
  assign k_sva_1_mx2_3 = MUX_s_1_2_2((k_sva_1[3]), (z_out_5_31_0[3]), fsm_output[13]);
  assign loop_1_loop_1_nand_seb_1 = ~((k_sva_1_mx1[7:6]==2'b11) & k_sva_1_mx2_3 &
      (~((k_sva_1_mx1[31]) | (k_sva_1_mx1[30]) | (k_sva_1_mx1[29]) | (k_sva_1_mx1[28])
      | (k_sva_1_mx1[27]) | (k_sva_1_mx1[26]) | (k_sva_1_mx1[25]) | (k_sva_1_mx1[24])
      | (k_sva_1_mx1[23]) | (k_sva_1_mx1[22]) | (k_sva_1_mx1[21]) | (k_sva_1_mx1[20])
      | (k_sva_1_mx1[19]) | (k_sva_1_mx1[18]) | (k_sva_1_mx1[17]) | (k_sva_1_mx1[16])
      | (k_sva_1_mx1[15]) | (k_sva_1_mx1[14]) | (k_sva_1_mx1[13]) | (k_sva_1_mx1[12])
      | (k_sva_1_mx1[11]) | (k_sva_1_mx1[10]) | (k_sva_1_mx1[9]) | (k_sva_1_mx1[8])
      | (k_sva_1_mx1[5]) | (k_sva_1_mx1[4]) | (k_sva_1_mx1[2]) | (k_sva_1_mx1[1])
      | (k_sva_1_mx1[0]))));
  assign and_dcpl_49 = ~((fsm_output[16]) | (fsm_output[17]) | (fsm_output[13]));
  assign or_dcpl_81 = (fsm_output[17]) | (fsm_output[13]);
  assign or_dcpl_83 = (fsm_output[15:14]!=2'b00);
  assign or_dcpl_85 = (fsm_output[18]) | (fsm_output[16]);
  assign or_tmp_46 = (fsm_output[10]) | (fsm_output[3]);
  assign j_3_0_sva_mx0c1 = (fsm_output[12]) | (fsm_output[17]) | ((z_out_3[4]) &
      (fsm_output[6]));
  assign j_3_0_sva_mx0c2 = (fsm_output[2]) | (fsm_output[13]) | ((~ loop_3_slc_loop_3_acc_3_itm)
      & (fsm_output[9])) | ((~ (z_out_3[4])) & (fsm_output[6]));
  assign row_buf_rsci_radr_d = row_buf_rsci_radr_d_reg;
  assign row_buf_rsci_wadr_d = row_buf_rsci_wadr_d_reg;
  assign row_buf_rsci_d_d = row_buf_rsci_d_d_reg;
  assign row_buf_rsci_we_d = row_buf_rsci_we_d_reg;
  assign row_buf_rsci_re_d = row_buf_rsci_re_d_reg;
  assign win_buf_rsci_radr_d = win_buf_rsci_radr_d_reg;
  assign win_buf_rsci_wadr_d = win_buf_rsci_wadr_d_reg;
  assign win_buf_rsci_d_d = win_buf_rsci_d_d_reg;
  assign win_buf_rsci_we_d = win_buf_rsci_we_d_reg;
  assign win_buf_rsci_re_d = win_buf_rsci_re_d_reg;
  assign or_tmp_86 = (fsm_output[17]) | (fsm_output[6]);
  assign or_tmp_89 = (fsm_output[17]) | (fsm_output[6]) | (fsm_output[12]) | (fsm_output[7]);
  assign loop_1_or_3_ssc = or_tmp_89 | (fsm_output[3]) | (fsm_output[14]);
  assign loop_8_or_ssc = or_tmp_46 | (fsm_output[13]);
  always @(posedge clk) begin
    if ( and_cse ) begin
      loop_op_i_15_0_sva <= loop_1_loop_1_and_2_cse;
      i_15_0_sva <= MUX_v_16_2_2(16'b0000000000000000, i_15_0_sva_2, (not_111_nl));
    end
  end
  always @(posedge clk) begin
    if ( core_wen & (fsm_output[18]) ) begin
      OUTPUT_rsci_idat_0 <= z_out_4[32];
    end
  end
  always @(posedge clk) begin
    if ( core_wen & ((fsm_output[0]) | (fsm_output[16]) | (fsm_output[17]) | (fsm_output[13])
        | (fsm_output[14]) | (fsm_output[19])) ) begin
      k_sva_31_8 <= MUX_v_24_2_2(24'b000000000000000000000000, (k_mux_5_nl), (k_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( core_wen ) begin
      k_sva_7_6 <= MUX_v_2_2_2(2'b00, (k_mux_4_nl), (nor_37_nl));
      k_sva_3 <= (k_mux1h_10_nl) & (~((fsm_output[16]) | (fsm_output[0])));
      loop_8_acc_10_itm <= MUX_v_6_2_2(z_out_7, ({3'b000 , (k_k_and_nl)}), nor_31_nl);
      loop_1_z_3_0_sva <= MUX_v_4_2_2(4'b0000, (n_mux1h_nl), (nor_nl));
      loop_3_acc_14_psp <= z_out;
      loop_3_acc_12_sdt_3_0 <= z_out_2_3_0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_INPUT_rsci_oswt_cse <= 1'b0;
      reg_OUTPUT_rsci_oswt_cse <= 1'b0;
      reg_row_buf_rsci_oswt_cse <= 1'b0;
      reg_win_buf_rsci_oswt_cse <= 1'b0;
      loop_lmm_loop_lmm_nor_itm <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_INPUT_rsci_oswt_cse <= ~((~((fsm_output[19]) | (fsm_output[0]))) | (loop_lmm_loop_lmm_nor_itm
          & (fsm_output[19])));
      reg_OUTPUT_rsci_oswt_cse <= fsm_output[18];
      reg_row_buf_rsci_oswt_cse <= or_141_rmff;
      reg_win_buf_rsci_oswt_cse <= or_tmp_46;
      loop_lmm_loop_lmm_nor_itm <= ~((readslicef_11_1_10((loop_lmm_acc_nl))) | (z_out_5_31_0[10])
          | (readslicef_11_1_10((loop_op_acc_nl))));
    end
  end
  always @(posedge clk) begin
    if ( core_wen & ((fsm_output[0]) | (fsm_output[19])) ) begin
      k_sva_5_4 <= MUX_v_2_2_2(2'b00, (k_sva_1[5:4]), (fsm_output[19]));
    end
  end
  always @(posedge clk) begin
    if ( ((fsm_output[1:0]!=2'b00)) & core_wen ) begin
      loop_lmm_i_15_0_sva <= loop_1_loop_1_and_2_cse;
    end
  end
  always @(posedge clk) begin
    if ( core_wen & ((loop_3_slc_loop_3_acc_3_itm & (fsm_output[9])) | j_3_0_sva_mx0c1
        | j_3_0_sva_mx0c2) ) begin
      j_3_0_sva <= MUX_v_4_2_2(4'b0000, (loop_1_z_mux_nl), (j_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( core_wen & ((fsm_output[7]) | or_tmp_46) ) begin
      loop_3_slc_loop_3_acc_3_itm <= z_out_1_3;
    end
  end
  always @(posedge clk) begin
    if ( core_wen & ((fsm_output[11]) | (fsm_output[9])) ) begin
      loop_1_sad_lpi_4 <= MUX_v_32_2_2(32'b00000000000000000000000000000000, (z_out_4[31:0]),
          (fsm_output[11]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      k_sva_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_85 | (fsm_output[17]) | or_dcpl_83)) ) begin
      k_sva_1 <= z_out_5_31_0;
    end
  end
  always @(posedge clk) begin
    if ( core_wen & (fsm_output[14]) ) begin
      o_7_0_sva_1 <= z_out_3;
    end
  end
  assign not_111_nl = ~ (fsm_output[0]);
  assign loop_8_mux_1_nl = MUX_v_8_2_2((k_sva_31_8[7:0]), o_7_0_sva_1, fsm_output[16]);
  assign or_211_nl = (fsm_output[16]) | (fsm_output[14]);
  assign loop_8_loop_8_and_nl = MUX_v_8_2_2(8'b00000000, (loop_8_mux_1_nl), (or_211_nl));
  assign k_mux_5_nl = MUX_v_24_2_2(({16'b0000000000000000 , (loop_8_loop_8_and_nl)}),
      (k_sva_1[31:8]), fsm_output[19]);
  assign k_not_nl = ~ (fsm_output[0]);
  assign nor_29_nl = ~((~ and_dcpl_49) | (fsm_output[14]) | (fsm_output[15]) | (fsm_output[0]));
  assign k_mux_4_nl = MUX_v_2_2_2((k_sva_1_mx1[7:6]), k_sva_7_6, nor_29_nl);
  assign nor_37_nl = ~((fsm_output[0]) | (fsm_output[14]) | (fsm_output[15]) | (fsm_output[16])
      | (~(and_dcpl_49 | loop_1_loop_1_nand_seb_1)));
  assign loop_1_loop_1_and_nl = k_sva_1_mx2_3 & loop_1_loop_1_nand_seb_1;
  assign and_146_nl = and_dcpl_49 & (~ (fsm_output[14])) & (~ (fsm_output[0]));
  assign k_mux1h_10_nl = MUX1HOT_s_1_3_2((loop_1_loop_1_and_nl), (z_out_5_31_0[5]),
      k_sva_3, {or_dcpl_81 , (fsm_output[14]) , (and_146_nl)});
  assign k_mux_3_nl = MUX_v_3_2_2((loop_8_acc_10_itm[2:0]), (k_sva_1[2:0]), fsm_output[19]);
  assign nor_32_nl = ~(or_dcpl_85 | or_dcpl_81 | or_dcpl_83 | (fsm_output[0]));
  assign k_k_and_nl = MUX_v_3_2_2(3'b000, (k_mux_3_nl), (nor_32_nl));
  assign nor_31_nl = ~((fsm_output[18:13]!=6'b000000));
  assign or_163_nl = (fsm_output[8]) | (fsm_output[5]) | (fsm_output[11]) | (fsm_output[4]);
  assign n_mux1h_nl = MUX1HOT_v_4_3_2((z_out_5_31_0[3:0]), loop_1_z_3_0_sva, (z_out_4[3:0]),
      {or_tmp_46 , (or_163_nl) , (fsm_output[7])});
  assign nor_nl = ~((fsm_output[2]) | (fsm_output[6]) | (fsm_output[12]) | (fsm_output[9]));
  assign nl_loop_lmm_acc_nl = conv_u2s_10_11(loop_lmm_i_15_0_sva[15:6]) + 11'b10110001111;
  assign loop_lmm_acc_nl = nl_loop_lmm_acc_nl[10:0];
  assign nl_loop_op_acc_nl = conv_u2s_10_11(z_out_6[15:6]) + 11'b10110001111;
  assign loop_op_acc_nl = nl_loop_op_acc_nl[10:0];
  assign loop_1_z_mux_nl = MUX_v_4_2_2(loop_1_z_3_0_sva, (z_out_4[3:0]), j_3_0_sva_mx0c1);
  assign j_not_nl = ~ j_3_0_sva_mx0c2;
  assign loop_3_or_4_nl = or_141_rmff | (fsm_output[10]);
  assign loop_3_mux_5_nl = MUX_v_4_2_2(loop_1_z_3_0_sva, j_3_0_sva, loop_3_or_4_nl);
  assign loop_3_loop_3_mux_1_nl = MUX_v_2_2_2((z_out_2_3_0[3:2]), (j_3_0_sva[3:2]),
      or_141_rmff);
  assign nl_z_out = (loop_3_mux_5_nl) + conv_u2u_2_4(loop_3_loop_3_mux_1_nl);
  assign z_out = nl_z_out[3:0];
  assign or_218_ssc = (fsm_output[12]) | (fsm_output[7]);
  assign loop_3_mux_6_nl = MUX_s_1_2_2((z_out_5_31_0[1]), (z_out_4[1]), or_218_ssc);
  assign loop_3_mux_7_nl = MUX_s_1_2_2((z_out_5_31_0[2]), (z_out_4[2]), or_218_ssc);
  assign loop_3_mux_8_nl = MUX_s_1_2_2((z_out_5_31_0[3]), (z_out_4[3]), or_218_ssc);
  assign z_out_1_3 = ~(((loop_3_mux_6_nl) | (loop_3_mux_7_nl)) & (loop_3_mux_8_nl));
  assign loop_4_mux_1_nl = MUX_v_4_2_2(j_3_0_sva, loop_1_z_3_0_sva, fsm_output[3]);
  assign loop_4_or_1_nl = (~((fsm_output[3]) | (fsm_output[10]))) | (fsm_output[7]);
  assign loop_4_mux1h_1_nl = MUX1HOT_v_3_3_2(({1'b0 , (j_3_0_sva[3:2])}), (j_3_0_sva[3:1]),
      (loop_1_z_3_0_sva[3:1]), {(fsm_output[7]) , (fsm_output[3]) , (fsm_output[10])});
  assign nl_acc_2_nl = ({(loop_4_mux_1_nl) , (loop_4_or_1_nl)}) + conv_u2u_4_5({(loop_4_mux1h_1_nl)
      , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[4:0];
  assign z_out_2_3_0 = readslicef_5_4_1((acc_2_nl));
  assign loop_8_mux_7_nl = MUX_v_8_2_2((k_sva_31_8[7:0]), 8'b11110111, or_tmp_86);
  assign loop_8_mux_8_nl = MUX_v_4_2_2(4'b0001, (z_out_4[3:0]), or_tmp_86);
  assign nl_z_out_3 = (loop_8_mux_7_nl) + conv_u2u_4_8(loop_8_mux_8_nl);
  assign z_out_3 = nl_z_out_3[7:0];
  assign loop_1_or_4_nl = (fsm_output[18]) | (fsm_output[11]);
  assign loop_1_or_5_nl = or_tmp_89 | (fsm_output[3]);
  assign loop_1_mux1h_4_nl = MUX1HOT_v_32_4_2(loop_1_sad_lpi_4, ({{28{j_3_0_sva[3]}},
      j_3_0_sva}), ({30'b000000000000000000000000000000 , (j_3_0_sva[3:2])}), (signext_32_6({(k_sva_7_6[0])
      , k_sva_5_4 , k_sva_3 , (loop_8_acc_10_itm[2:1])})), {(loop_1_or_4_nl) , (loop_1_or_5_nl)
      , (fsm_output[14]) , (fsm_output[1])});
  assign loop_1_loop_1_or_1_nl = (~((fsm_output[11]) | loop_1_or_3_ssc)) | (fsm_output[1]);
  assign loop_1_mux1h_5_nl = MUX1HOT_v_8_3_2(win_buf_rsci_q_d_mxwt, 8'b00000001,
      8'b11101101, {(fsm_output[11]) , loop_1_or_3_ssc , (fsm_output[1])});
  assign loop_1_or_6_nl = MUX_v_9_2_2(({(loop_1_loop_1_or_1_nl) , (loop_1_mux1h_5_nl)}),
      9'b111111111, (fsm_output[18]));
  assign nl_z_out_4 = conv_s2u_32_33(loop_1_mux1h_4_nl) + conv_s2u_9_33(loop_1_or_6_nl);
  assign z_out_4 = nl_z_out_4[32:0];
  assign loop_8_mux1h_4_nl = MUX1HOT_v_32_4_2(({27'b000000000000000000000000000 ,
      (z_out_3[7:3])}), ({{28{loop_1_z_3_0_sva[3]}}, loop_1_z_3_0_sva}), ({k_sva_31_8
      , k_sva_7_6 , k_sva_5_4 , k_sva_3 , (loop_8_acc_10_itm[2:0])}), ({22'b0000000000000000000000
      , (i_15_0_sva_2[15:6])}), {(fsm_output[14]) , or_tmp_46 , (fsm_output[13])
      , (fsm_output[18])});
  assign loop_8_loop_8_or_3_nl = (~ loop_8_or_ssc) | (fsm_output[14]);
  assign loop_8_not_4_nl = ~ loop_8_or_ssc;
  assign loop_8_loop_8_or_4_nl = MUX_v_2_2_2((signext_2_1(fsm_output[14])), 2'b11,
      (loop_8_not_4_nl));
  assign loop_8_not_5_nl = ~ loop_8_or_ssc;
  assign loop_8_loop_8_or_5_nl = MUX_v_2_2_2((signext_2_1(fsm_output[18])), 2'b11,
      (loop_8_not_5_nl));
  assign nl_z_out_5_31_0 = (loop_8_mux1h_4_nl) + conv_s2u_11_32({(loop_8_loop_8_or_3_nl)
      , (fsm_output[14]) , (loop_8_loop_8_or_4_nl) , (signext_2_1(fsm_output[14]))
      , 1'b0 , (fsm_output[18]) , (loop_8_loop_8_or_5_nl) , 1'b1});
  assign z_out_5_31_0 = nl_z_out_5_31_0[31:0];
  assign loop_lmm_mux_3_nl = MUX_v_16_2_2(loop_lmm_i_15_0_sva, loop_op_i_15_0_sva,
      fsm_output[18]);
  assign nl_z_out_6 = (loop_lmm_mux_3_nl) + 16'b0000000000000001;
  assign z_out_6 = nl_z_out_6[15:0];
  assign loop_8_mux_9_nl = MUX_v_6_2_2((k_sva_31_8[6:1]), ({(k_sva_7_6[0]) , k_sva_5_4
      , k_sva_3 , (loop_8_acc_10_itm[2:1])}), fsm_output[7]);
  assign nl_z_out_7 = ({z_out , (j_3_0_sva[1:0])}) + (loop_8_mux_9_nl);
  assign z_out_7 = nl_z_out_7[5:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_4_2;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [3:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    MUX1HOT_v_32_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [23:0] MUX_v_24_2_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input [0:0] sel;
    reg [23:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_24_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [3:0] readslicef_5_4_1;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_5_4_1 = tmp[3:0];
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [31:0] signext_32_6;
    input [5:0] vector;
  begin
    signext_32_6= {{26{vector[5]}}, vector};
  end
  endfunction


  function automatic [32:0] conv_s2u_9_33 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_33 = {{24{vector[8]}}, vector};
  end
  endfunction


  function automatic [31:0] conv_s2u_11_32 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_32 = {{21{vector[10]}}, vector};
  end
  endfunction


  function automatic [32:0] conv_s2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_s2u_32_33 = {vector[31], vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_4_6 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_6 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_4_8 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_8 = {{4{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SAD_MATCH
// ------------------------------------------------------------------


module SAD_MATCH (
  clk, rst, INPUT_rsc_dat, INPUT_rsc_vld, INPUT_rsc_rdy, OUTPUT_rsc_dat, OUTPUT_rsc_vld,
      OUTPUT_rsc_rdy
);
  input clk;
  input rst;
  input [7:0] INPUT_rsc_dat;
  input INPUT_rsc_vld;
  output INPUT_rsc_rdy;
  output [7:0] OUTPUT_rsc_dat;
  output OUTPUT_rsc_vld;
  input OUTPUT_rsc_rdy;


  // Interconnect Declarations
  wire [6:0] row_buf_rsci_radr_d;
  wire [6:0] row_buf_rsci_wadr_d;
  wire [7:0] row_buf_rsci_d_d;
  wire row_buf_rsci_we_d;
  wire row_buf_rsci_re_d;
  wire [7:0] row_buf_rsci_q_d;
  wire [6:0] win_buf_rsci_radr_d;
  wire [6:0] win_buf_rsci_wadr_d;
  wire [7:0] win_buf_rsci_d_d;
  wire win_buf_rsci_we_d;
  wire win_buf_rsci_re_d;
  wire [7:0] win_buf_rsci_q_d;
  wire row_buf_rsc_we;
  wire [7:0] row_buf_rsc_d;
  wire [6:0] row_buf_rsc_wadr;
  wire row_buf_rsc_re;
  wire [7:0] row_buf_rsc_q;
  wire [6:0] row_buf_rsc_radr;
  wire win_buf_rsc_we;
  wire [7:0] win_buf_rsc_d;
  wire [6:0] win_buf_rsc_wadr;
  wire win_buf_rsc_re;
  wire [7:0] win_buf_rsc_q;
  wire [6:0] win_buf_rsc_radr;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.data_width(32'sd8),
  .addr_width(32'sd7),
  .depth(32'sd100)) row_buf_rsc_comp (
      .radr(row_buf_rsc_radr),
      .wadr(row_buf_rsc_wadr),
      .d(row_buf_rsc_d),
      .we(row_buf_rsc_we),
      .re(row_buf_rsc_re),
      .clk(clk),
      .q(row_buf_rsc_q)
    );
  BLOCK_1R1W_RBW #(.data_width(32'sd8),
  .addr_width(32'sd7),
  .depth(32'sd100)) win_buf_rsc_comp (
      .radr(win_buf_rsc_radr),
      .wadr(win_buf_rsc_wadr),
      .d(win_buf_rsc_d),
      .we(win_buf_rsc_we),
      .re(win_buf_rsc_re),
      .clk(clk),
      .q(win_buf_rsc_q)
    );
  SAD_MATCH_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_7_100_5_gen row_buf_rsci (
      .we(row_buf_rsc_we),
      .d(row_buf_rsc_d),
      .wadr(row_buf_rsc_wadr),
      .re(row_buf_rsc_re),
      .q(row_buf_rsc_q),
      .radr(row_buf_rsc_radr),
      .radr_d(row_buf_rsci_radr_d),
      .wadr_d(row_buf_rsci_wadr_d),
      .d_d(row_buf_rsci_d_d),
      .we_d(row_buf_rsci_we_d),
      .re_d(row_buf_rsci_re_d),
      .q_d(row_buf_rsci_q_d)
    );
  SAD_MATCH_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_7_100_6_gen win_buf_rsci (
      .we(win_buf_rsc_we),
      .d(win_buf_rsc_d),
      .wadr(win_buf_rsc_wadr),
      .re(win_buf_rsc_re),
      .q(win_buf_rsc_q),
      .radr(win_buf_rsc_radr),
      .radr_d(win_buf_rsci_radr_d),
      .wadr_d(win_buf_rsci_wadr_d),
      .d_d(win_buf_rsci_d_d),
      .we_d(win_buf_rsci_we_d),
      .re_d(win_buf_rsci_re_d),
      .q_d(win_buf_rsci_q_d)
    );
  SAD_MATCH_core SAD_MATCH_core_inst (
      .clk(clk),
      .rst(rst),
      .INPUT_rsc_dat(INPUT_rsc_dat),
      .INPUT_rsc_vld(INPUT_rsc_vld),
      .INPUT_rsc_rdy(INPUT_rsc_rdy),
      .OUTPUT_rsc_dat(OUTPUT_rsc_dat),
      .OUTPUT_rsc_vld(OUTPUT_rsc_vld),
      .OUTPUT_rsc_rdy(OUTPUT_rsc_rdy),
      .row_buf_rsci_radr_d(row_buf_rsci_radr_d),
      .row_buf_rsci_wadr_d(row_buf_rsci_wadr_d),
      .row_buf_rsci_d_d(row_buf_rsci_d_d),
      .row_buf_rsci_we_d(row_buf_rsci_we_d),
      .row_buf_rsci_re_d(row_buf_rsci_re_d),
      .row_buf_rsci_q_d(row_buf_rsci_q_d),
      .win_buf_rsci_radr_d(win_buf_rsci_radr_d),
      .win_buf_rsci_wadr_d(win_buf_rsci_wadr_d),
      .win_buf_rsci_d_d(win_buf_rsci_d_d),
      .win_buf_rsci_we_d(win_buf_rsci_we_d),
      .win_buf_rsci_re_d(win_buf_rsci_re_d),
      .win_buf_rsci_q_d(win_buf_rsci_q_d)
    );
endmodule



