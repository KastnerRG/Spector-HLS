
//------> /usr/local/bin/Mentor_Graphics/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /usr/local/bin/Mentor_Graphics/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /usr/local/bin/Mentor_Graphics/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Block 1R1W Read Before Write RAM with common clock
module BLOCK_1R1W_RBW
#(
parameter data_width = 8,
parameter addr_width = 7,
parameter depth = 128
)(
	radr, wadr, d, we, re, clk, q
);

	input [addr_width-1:0] radr;
	input [addr_width-1:0] wadr;
	input [data_width-1:0] d;
	input we;
	input re;
	input clk;
	output[data_width-1:0] q;

	reg [data_width-1:0] q;

	(* ram_style = "block" *)
	reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block_ram"
	//pragma attribute mem block_ram true
		
	always @(posedge clk) begin
		if (we) begin
			mem[wadr] <= d; // Write port
		end
		if (re) begin
			q <= mem[radr] ; // read port
		end
	end

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   mdk@mdk-FX504
//  Generated date: Fri Feb 14 16:11:01 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    DCT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_22_4194304_4_gen
// ------------------------------------------------------------------


module DCT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_22_4194304_4_gen (
  we, d, wadr, re, q, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d
);
  output we;
  output [19:0] d;
  output [21:0] wadr;
  output re;
  input [19:0] q;
  output [21:0] radr;
  input [21:0] radr_d;
  input [21:0] wadr_d;
  input [19:0] d_d;
  input we_d;
  input re_d;
  output [19:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_22_4194304_3_gen
// ------------------------------------------------------------------


module DCT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_22_4194304_3_gen (
  we, d, wadr, re, q, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d
);
  output we;
  output [19:0] d;
  output [21:0] wadr;
  output re;
  input [19:0] q;
  output [21:0] radr;
  input [21:0] radr_d;
  input [21:0] wadr_d;
  input [19:0] d_d;
  input we_d;
  input re_d;
  output [19:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module DCT_core_core_fsm (
  clk, rst, core_wen, fsm_output, loop_lmm_C_1_tr0, loop_6_C_2_tr0, loop_5_C_1_tr0,
      loop_7_C_1_tr0, loop_7_C_1_tr1, loop_3_C_0_tr0, loop_12_C_2_tr0, loop_11_C_1_tr0,
      loop_13_C_1_tr0, loop_13_C_1_tr1, loop_9_C_0_tr0, loop_2_C_0_tr0, loop_1_C_0_tr0,
      loop_out_C_2_tr0
);
  input clk;
  input rst;
  input core_wen;
  output [27:0] fsm_output;
  reg [27:0] fsm_output;
  input loop_lmm_C_1_tr0;
  input loop_6_C_2_tr0;
  input loop_5_C_1_tr0;
  input loop_7_C_1_tr0;
  input loop_7_C_1_tr1;
  input loop_3_C_0_tr0;
  input loop_12_C_2_tr0;
  input loop_11_C_1_tr0;
  input loop_13_C_1_tr0;
  input loop_13_C_1_tr1;
  input loop_9_C_0_tr0;
  input loop_2_C_0_tr0;
  input loop_1_C_0_tr0;
  input loop_out_C_2_tr0;


  // FSM State Type Declaration for DCT_core_core_fsm_1
  parameter
    main_C_0 = 5'd0,
    loop_lmm_C_0 = 5'd1,
    loop_lmm_C_1 = 5'd2,
    loop_5_C_0 = 5'd3,
    loop_6_C_0 = 5'd4,
    loop_6_C_1 = 5'd5,
    loop_6_C_2 = 5'd6,
    loop_5_C_1 = 5'd7,
    loop_4_C_0 = 5'd8,
    loop_4_C_1 = 5'd9,
    loop_7_C_0 = 5'd10,
    loop_7_C_1 = 5'd11,
    loop_3_C_0 = 5'd12,
    loop_11_C_0 = 5'd13,
    loop_12_C_0 = 5'd14,
    loop_12_C_1 = 5'd15,
    loop_12_C_2 = 5'd16,
    loop_11_C_1 = 5'd17,
    loop_10_C_0 = 5'd18,
    loop_10_C_1 = 5'd19,
    loop_13_C_0 = 5'd20,
    loop_13_C_1 = 5'd21,
    loop_9_C_0 = 5'd22,
    loop_2_C_0 = 5'd23,
    loop_1_C_0 = 5'd24,
    loop_out_C_0 = 5'd25,
    loop_out_C_1 = 5'd26,
    loop_out_C_2 = 5'd27;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : DCT_core_core_fsm_1
    case (state_var)
      loop_lmm_C_0 : begin
        fsm_output = 28'b0000000000000000000000000010;
        state_var_NS = loop_lmm_C_1;
      end
      loop_lmm_C_1 : begin
        fsm_output = 28'b0000000000000000000000000100;
        if ( loop_lmm_C_1_tr0 ) begin
          state_var_NS = loop_5_C_0;
        end
        else begin
          state_var_NS = loop_lmm_C_0;
        end
      end
      loop_5_C_0 : begin
        fsm_output = 28'b0000000000000000000000001000;
        state_var_NS = loop_6_C_0;
      end
      loop_6_C_0 : begin
        fsm_output = 28'b0000000000000000000000010000;
        state_var_NS = loop_6_C_1;
      end
      loop_6_C_1 : begin
        fsm_output = 28'b0000000000000000000000100000;
        state_var_NS = loop_6_C_2;
      end
      loop_6_C_2 : begin
        fsm_output = 28'b0000000000000000000001000000;
        if ( loop_6_C_2_tr0 ) begin
          state_var_NS = loop_5_C_1;
        end
        else begin
          state_var_NS = loop_6_C_0;
        end
      end
      loop_5_C_1 : begin
        fsm_output = 28'b0000000000000000000010000000;
        if ( loop_5_C_1_tr0 ) begin
          state_var_NS = loop_4_C_0;
        end
        else begin
          state_var_NS = loop_5_C_0;
        end
      end
      loop_4_C_0 : begin
        fsm_output = 28'b0000000000000000000100000000;
        state_var_NS = loop_4_C_1;
      end
      loop_4_C_1 : begin
        fsm_output = 28'b0000000000000000001000000000;
        state_var_NS = loop_7_C_0;
      end
      loop_7_C_0 : begin
        fsm_output = 28'b0000000000000000010000000000;
        state_var_NS = loop_7_C_1;
      end
      loop_7_C_1 : begin
        fsm_output = 28'b0000000000000000100000000000;
        if ( loop_7_C_1_tr0 ) begin
          state_var_NS = loop_3_C_0;
        end
        else if ( loop_7_C_1_tr1 ) begin
          state_var_NS = loop_7_C_0;
        end
        else begin
          state_var_NS = loop_5_C_0;
        end
      end
      loop_3_C_0 : begin
        fsm_output = 28'b0000000000000001000000000000;
        if ( loop_3_C_0_tr0 ) begin
          state_var_NS = loop_11_C_0;
        end
        else begin
          state_var_NS = loop_5_C_0;
        end
      end
      loop_11_C_0 : begin
        fsm_output = 28'b0000000000000010000000000000;
        state_var_NS = loop_12_C_0;
      end
      loop_12_C_0 : begin
        fsm_output = 28'b0000000000000100000000000000;
        state_var_NS = loop_12_C_1;
      end
      loop_12_C_1 : begin
        fsm_output = 28'b0000000000001000000000000000;
        state_var_NS = loop_12_C_2;
      end
      loop_12_C_2 : begin
        fsm_output = 28'b0000000000010000000000000000;
        if ( loop_12_C_2_tr0 ) begin
          state_var_NS = loop_11_C_1;
        end
        else begin
          state_var_NS = loop_12_C_0;
        end
      end
      loop_11_C_1 : begin
        fsm_output = 28'b0000000000100000000000000000;
        if ( loop_11_C_1_tr0 ) begin
          state_var_NS = loop_10_C_0;
        end
        else begin
          state_var_NS = loop_11_C_0;
        end
      end
      loop_10_C_0 : begin
        fsm_output = 28'b0000000001000000000000000000;
        state_var_NS = loop_10_C_1;
      end
      loop_10_C_1 : begin
        fsm_output = 28'b0000000010000000000000000000;
        state_var_NS = loop_13_C_0;
      end
      loop_13_C_0 : begin
        fsm_output = 28'b0000000100000000000000000000;
        state_var_NS = loop_13_C_1;
      end
      loop_13_C_1 : begin
        fsm_output = 28'b0000001000000000000000000000;
        if ( loop_13_C_1_tr0 ) begin
          state_var_NS = loop_9_C_0;
        end
        else if ( loop_13_C_1_tr1 ) begin
          state_var_NS = loop_13_C_0;
        end
        else begin
          state_var_NS = loop_11_C_0;
        end
      end
      loop_9_C_0 : begin
        fsm_output = 28'b0000010000000000000000000000;
        if ( loop_9_C_0_tr0 ) begin
          state_var_NS = loop_2_C_0;
        end
        else begin
          state_var_NS = loop_11_C_0;
        end
      end
      loop_2_C_0 : begin
        fsm_output = 28'b0000100000000000000000000000;
        if ( loop_2_C_0_tr0 ) begin
          state_var_NS = loop_1_C_0;
        end
        else begin
          state_var_NS = loop_5_C_0;
        end
      end
      loop_1_C_0 : begin
        fsm_output = 28'b0001000000000000000000000000;
        if ( loop_1_C_0_tr0 ) begin
          state_var_NS = loop_out_C_0;
        end
        else begin
          state_var_NS = loop_5_C_0;
        end
      end
      loop_out_C_0 : begin
        fsm_output = 28'b0010000000000000000000000000;
        state_var_NS = loop_out_C_1;
      end
      loop_out_C_1 : begin
        fsm_output = 28'b0100000000000000000000000000;
        state_var_NS = loop_out_C_2;
      end
      loop_out_C_2 : begin
        fsm_output = 28'b1000000000000000000000000000;
        if ( loop_out_C_2_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = loop_out_C_0;
        end
      end
      // main_C_0
      default : begin
        fsm_output = 28'b0000000000000000000000000001;
        state_var_NS = loop_lmm_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_staller
// ------------------------------------------------------------------


module DCT_core_staller (
  clk, rst, core_wen, core_wten, dst_rsci_wen_comp, src_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input dst_rsci_wen_comp;
  input src_rsci_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = dst_rsci_wen_comp & src_rsci_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_msrc_data_rsci_1_msrc_data_rsc_wait_dp
// ------------------------------------------------------------------


module DCT_core_msrc_data_rsci_1_msrc_data_rsc_wait_dp (
  clk, rst, msrc_data_rsci_radr_d, msrc_data_rsci_wadr_d, msrc_data_rsci_d_d, msrc_data_rsci_q_d,
      msrc_data_rsci_radr_d_core, msrc_data_rsci_wadr_d_core, msrc_data_rsci_d_d_core,
      msrc_data_rsci_q_d_mxwt, msrc_data_rsci_biwt, msrc_data_rsci_bdwt, msrc_data_rsci_radr_d_core_sct,
      msrc_data_rsci_wadr_d_core_sct_pff
);
  input clk;
  input rst;
  output [21:0] msrc_data_rsci_radr_d;
  output [21:0] msrc_data_rsci_wadr_d;
  output [19:0] msrc_data_rsci_d_d;
  input [19:0] msrc_data_rsci_q_d;
  input [21:0] msrc_data_rsci_radr_d_core;
  input [21:0] msrc_data_rsci_wadr_d_core;
  input [19:0] msrc_data_rsci_d_d_core;
  output [19:0] msrc_data_rsci_q_d_mxwt;
  input msrc_data_rsci_biwt;
  input msrc_data_rsci_bdwt;
  input msrc_data_rsci_radr_d_core_sct;
  input msrc_data_rsci_wadr_d_core_sct_pff;


  // Interconnect Declarations
  reg msrc_data_rsci_bcwt;
  reg [19:0] msrc_data_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign msrc_data_rsci_q_d_mxwt = MUX_v_20_2_2(msrc_data_rsci_q_d, msrc_data_rsci_q_d_bfwt,
      msrc_data_rsci_bcwt);
  assign msrc_data_rsci_radr_d = MUX_v_22_2_2(22'b0000000000000000000000, msrc_data_rsci_radr_d_core,
      msrc_data_rsci_radr_d_core_sct);
  assign msrc_data_rsci_wadr_d = MUX_v_22_2_2(22'b0000000000000000000000, msrc_data_rsci_wadr_d_core,
      msrc_data_rsci_wadr_d_core_sct_pff);
  assign msrc_data_rsci_d_d = MUX_v_20_2_2(20'b00000000000000000000, msrc_data_rsci_d_d_core,
      msrc_data_rsci_wadr_d_core_sct_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      msrc_data_rsci_bcwt <= 1'b0;
    end
    else begin
      msrc_data_rsci_bcwt <= ~((~(msrc_data_rsci_bcwt | msrc_data_rsci_biwt)) | msrc_data_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ msrc_data_rsci_bcwt ) begin
      msrc_data_rsci_q_d_bfwt <= msrc_data_rsci_q_d_mxwt;
    end
  end

  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_msrc_data_rsci_1_msrc_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module DCT_core_msrc_data_rsci_1_msrc_data_rsc_wait_ctrl (
  core_wen, core_wten, msrc_data_rsci_oswt, msrc_data_rsci_biwt, msrc_data_rsci_bdwt,
      msrc_data_rsci_radr_d_core_sct_pff, msrc_data_rsci_oswt_pff, msrc_data_rsci_wadr_d_core_sct_pff,
      msrc_data_rsci_iswt0_1_pff
);
  input core_wen;
  input core_wten;
  input msrc_data_rsci_oswt;
  output msrc_data_rsci_biwt;
  output msrc_data_rsci_bdwt;
  output msrc_data_rsci_radr_d_core_sct_pff;
  input msrc_data_rsci_oswt_pff;
  output msrc_data_rsci_wadr_d_core_sct_pff;
  input msrc_data_rsci_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign msrc_data_rsci_bdwt = msrc_data_rsci_oswt & core_wen;
  assign msrc_data_rsci_biwt = (~ core_wten) & msrc_data_rsci_oswt;
  assign msrc_data_rsci_radr_d_core_sct_pff = msrc_data_rsci_oswt_pff & core_wen;
  assign msrc_data_rsci_wadr_d_core_sct_pff = msrc_data_rsci_iswt0_1_pff & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_mdst_data_rsci_1_mdst_data_rsc_wait_dp
// ------------------------------------------------------------------


module DCT_core_mdst_data_rsci_1_mdst_data_rsc_wait_dp (
  clk, rst, mdst_data_rsci_radr_d, mdst_data_rsci_wadr_d, mdst_data_rsci_d_d, mdst_data_rsci_q_d,
      mdst_data_rsci_radr_d_core, mdst_data_rsci_wadr_d_core, mdst_data_rsci_d_d_core,
      mdst_data_rsci_q_d_mxwt, mdst_data_rsci_biwt, mdst_data_rsci_bdwt, mdst_data_rsci_radr_d_core_sct,
      mdst_data_rsci_wadr_d_core_sct_pff
);
  input clk;
  input rst;
  output [21:0] mdst_data_rsci_radr_d;
  output [21:0] mdst_data_rsci_wadr_d;
  output [19:0] mdst_data_rsci_d_d;
  input [19:0] mdst_data_rsci_q_d;
  input [21:0] mdst_data_rsci_radr_d_core;
  input [21:0] mdst_data_rsci_wadr_d_core;
  input [19:0] mdst_data_rsci_d_d_core;
  output [19:0] mdst_data_rsci_q_d_mxwt;
  input mdst_data_rsci_biwt;
  input mdst_data_rsci_bdwt;
  input mdst_data_rsci_radr_d_core_sct;
  input mdst_data_rsci_wadr_d_core_sct_pff;


  // Interconnect Declarations
  reg mdst_data_rsci_bcwt;
  reg [19:0] mdst_data_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign mdst_data_rsci_q_d_mxwt = MUX_v_20_2_2(mdst_data_rsci_q_d, mdst_data_rsci_q_d_bfwt,
      mdst_data_rsci_bcwt);
  assign mdst_data_rsci_radr_d = MUX_v_22_2_2(22'b0000000000000000000000, mdst_data_rsci_radr_d_core,
      mdst_data_rsci_radr_d_core_sct);
  assign mdst_data_rsci_wadr_d = MUX_v_22_2_2(22'b0000000000000000000000, mdst_data_rsci_wadr_d_core,
      mdst_data_rsci_wadr_d_core_sct_pff);
  assign mdst_data_rsci_d_d = MUX_v_20_2_2(20'b00000000000000000000, mdst_data_rsci_d_d_core,
      mdst_data_rsci_wadr_d_core_sct_pff);
  always @(posedge clk) begin
    if ( rst ) begin
      mdst_data_rsci_bcwt <= 1'b0;
    end
    else begin
      mdst_data_rsci_bcwt <= ~((~(mdst_data_rsci_bcwt | mdst_data_rsci_biwt)) | mdst_data_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ mdst_data_rsci_bcwt ) begin
      mdst_data_rsci_q_d_bfwt <= mdst_data_rsci_q_d_mxwt;
    end
  end

  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_mdst_data_rsci_1_mdst_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module DCT_core_mdst_data_rsci_1_mdst_data_rsc_wait_ctrl (
  core_wen, core_wten, mdst_data_rsci_oswt, mdst_data_rsci_biwt, mdst_data_rsci_bdwt,
      mdst_data_rsci_radr_d_core_sct_pff, mdst_data_rsci_oswt_pff, mdst_data_rsci_wadr_d_core_sct_pff,
      mdst_data_rsci_iswt0_1_pff
);
  input core_wen;
  input core_wten;
  input mdst_data_rsci_oswt;
  output mdst_data_rsci_biwt;
  output mdst_data_rsci_bdwt;
  output mdst_data_rsci_radr_d_core_sct_pff;
  input mdst_data_rsci_oswt_pff;
  output mdst_data_rsci_wadr_d_core_sct_pff;
  input mdst_data_rsci_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign mdst_data_rsci_bdwt = mdst_data_rsci_oswt & core_wen;
  assign mdst_data_rsci_biwt = (~ core_wten) & mdst_data_rsci_oswt;
  assign mdst_data_rsci_radr_d_core_sct_pff = mdst_data_rsci_oswt_pff & core_wen;
  assign mdst_data_rsci_wadr_d_core_sct_pff = mdst_data_rsci_iswt0_1_pff & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_src_rsci_src_wait_dp
// ------------------------------------------------------------------


module DCT_core_src_rsci_src_wait_dp (
  clk, rst, src_rsci_oswt, src_rsci_wen_comp, src_rsci_idat_mxwt, src_rsci_biwt,
      src_rsci_bdwt, src_rsci_bcwt, src_rsci_idat
);
  input clk;
  input rst;
  input src_rsci_oswt;
  output src_rsci_wen_comp;
  output [19:0] src_rsci_idat_mxwt;
  input src_rsci_biwt;
  input src_rsci_bdwt;
  output src_rsci_bcwt;
  reg src_rsci_bcwt;
  input [19:0] src_rsci_idat;


  // Interconnect Declarations
  reg [19:0] src_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign src_rsci_wen_comp = (~ src_rsci_oswt) | src_rsci_biwt | src_rsci_bcwt;
  assign src_rsci_idat_mxwt = MUX_v_20_2_2(src_rsci_idat, src_rsci_idat_bfwt, src_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      src_rsci_bcwt <= 1'b0;
    end
    else begin
      src_rsci_bcwt <= ~((~(src_rsci_bcwt | src_rsci_biwt)) | src_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    src_rsci_idat_bfwt <= src_rsci_idat_mxwt;
  end

  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_src_rsci_src_wait_ctrl
// ------------------------------------------------------------------


module DCT_core_src_rsci_src_wait_ctrl (
  core_wen, src_rsci_oswt, src_rsci_biwt, src_rsci_bdwt, src_rsci_bcwt, src_rsci_irdy_core_sct,
      src_rsci_ivld
);
  input core_wen;
  input src_rsci_oswt;
  output src_rsci_biwt;
  output src_rsci_bdwt;
  input src_rsci_bcwt;
  output src_rsci_irdy_core_sct;
  input src_rsci_ivld;


  // Interconnect Declarations
  wire src_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign src_rsci_bdwt = src_rsci_oswt & core_wen;
  assign src_rsci_biwt = src_rsci_ogwt & src_rsci_ivld;
  assign src_rsci_ogwt = src_rsci_oswt & (~ src_rsci_bcwt);
  assign src_rsci_irdy_core_sct = src_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_dst_rsci_dst_wait_dp
// ------------------------------------------------------------------


module DCT_core_dst_rsci_dst_wait_dp (
  clk, rst, dst_rsci_oswt, dst_rsci_wen_comp, dst_rsci_biwt, dst_rsci_bdwt, dst_rsci_bcwt
);
  input clk;
  input rst;
  input dst_rsci_oswt;
  output dst_rsci_wen_comp;
  input dst_rsci_biwt;
  input dst_rsci_bdwt;
  output dst_rsci_bcwt;
  reg dst_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dst_rsci_wen_comp = (~ dst_rsci_oswt) | dst_rsci_biwt | dst_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      dst_rsci_bcwt <= 1'b0;
    end
    else begin
      dst_rsci_bcwt <= ~((~(dst_rsci_bcwt | dst_rsci_biwt)) | dst_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_dst_rsci_dst_wait_ctrl
// ------------------------------------------------------------------


module DCT_core_dst_rsci_dst_wait_ctrl (
  core_wen, dst_rsci_oswt, dst_rsci_irdy, dst_rsci_biwt, dst_rsci_bdwt, dst_rsci_bcwt,
      dst_rsci_ivld_core_sct
);
  input core_wen;
  input dst_rsci_oswt;
  input dst_rsci_irdy;
  output dst_rsci_biwt;
  output dst_rsci_bdwt;
  input dst_rsci_bcwt;
  output dst_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire dst_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dst_rsci_bdwt = dst_rsci_oswt & core_wen;
  assign dst_rsci_biwt = dst_rsci_ogwt & dst_rsci_irdy;
  assign dst_rsci_ogwt = dst_rsci_oswt & (~ dst_rsci_bcwt);
  assign dst_rsci_ivld_core_sct = dst_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_msrc_data_rsci_1
// ------------------------------------------------------------------


module DCT_core_msrc_data_rsci_1 (
  clk, rst, msrc_data_rsci_radr_d, msrc_data_rsci_wadr_d, msrc_data_rsci_d_d, msrc_data_rsci_we_d,
      msrc_data_rsci_re_d, msrc_data_rsci_q_d, core_wen, core_wten, msrc_data_rsci_oswt,
      msrc_data_rsci_radr_d_core, msrc_data_rsci_wadr_d_core, msrc_data_rsci_d_d_core,
      msrc_data_rsci_q_d_mxwt, msrc_data_rsci_oswt_pff, msrc_data_rsci_iswt0_1_pff
);
  input clk;
  input rst;
  output [21:0] msrc_data_rsci_radr_d;
  output [21:0] msrc_data_rsci_wadr_d;
  output [19:0] msrc_data_rsci_d_d;
  output msrc_data_rsci_we_d;
  output msrc_data_rsci_re_d;
  input [19:0] msrc_data_rsci_q_d;
  input core_wen;
  input core_wten;
  input msrc_data_rsci_oswt;
  input [21:0] msrc_data_rsci_radr_d_core;
  input [21:0] msrc_data_rsci_wadr_d_core;
  input [19:0] msrc_data_rsci_d_d_core;
  output [19:0] msrc_data_rsci_q_d_mxwt;
  input msrc_data_rsci_oswt_pff;
  input msrc_data_rsci_iswt0_1_pff;


  // Interconnect Declarations
  wire msrc_data_rsci_biwt;
  wire msrc_data_rsci_bdwt;
  wire [21:0] msrc_data_rsci_radr_d_reg;
  wire msrc_data_rsci_radr_d_core_sct_iff;
  wire [21:0] msrc_data_rsci_wadr_d_reg;
  wire msrc_data_rsci_wadr_d_core_sct_iff;
  wire [19:0] msrc_data_rsci_d_d_reg;


  // Interconnect Declarations for Component Instantiations 
  DCT_core_msrc_data_rsci_1_msrc_data_rsc_wait_ctrl DCT_core_msrc_data_rsci_1_msrc_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .msrc_data_rsci_oswt(msrc_data_rsci_oswt),
      .msrc_data_rsci_biwt(msrc_data_rsci_biwt),
      .msrc_data_rsci_bdwt(msrc_data_rsci_bdwt),
      .msrc_data_rsci_radr_d_core_sct_pff(msrc_data_rsci_radr_d_core_sct_iff),
      .msrc_data_rsci_oswt_pff(msrc_data_rsci_oswt_pff),
      .msrc_data_rsci_wadr_d_core_sct_pff(msrc_data_rsci_wadr_d_core_sct_iff),
      .msrc_data_rsci_iswt0_1_pff(msrc_data_rsci_iswt0_1_pff)
    );
  DCT_core_msrc_data_rsci_1_msrc_data_rsc_wait_dp DCT_core_msrc_data_rsci_1_msrc_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .msrc_data_rsci_radr_d(msrc_data_rsci_radr_d_reg),
      .msrc_data_rsci_wadr_d(msrc_data_rsci_wadr_d_reg),
      .msrc_data_rsci_d_d(msrc_data_rsci_d_d_reg),
      .msrc_data_rsci_q_d(msrc_data_rsci_q_d),
      .msrc_data_rsci_radr_d_core(msrc_data_rsci_radr_d_core),
      .msrc_data_rsci_wadr_d_core(msrc_data_rsci_wadr_d_core),
      .msrc_data_rsci_d_d_core(msrc_data_rsci_d_d_core),
      .msrc_data_rsci_q_d_mxwt(msrc_data_rsci_q_d_mxwt),
      .msrc_data_rsci_biwt(msrc_data_rsci_biwt),
      .msrc_data_rsci_bdwt(msrc_data_rsci_bdwt),
      .msrc_data_rsci_radr_d_core_sct(msrc_data_rsci_radr_d_core_sct_iff),
      .msrc_data_rsci_wadr_d_core_sct_pff(msrc_data_rsci_wadr_d_core_sct_iff)
    );
  assign msrc_data_rsci_radr_d = msrc_data_rsci_radr_d_reg;
  assign msrc_data_rsci_wadr_d = msrc_data_rsci_wadr_d_reg;
  assign msrc_data_rsci_d_d = msrc_data_rsci_d_d_reg;
  assign msrc_data_rsci_we_d = msrc_data_rsci_wadr_d_core_sct_iff;
  assign msrc_data_rsci_re_d = msrc_data_rsci_radr_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_mdst_data_rsci_1
// ------------------------------------------------------------------


module DCT_core_mdst_data_rsci_1 (
  clk, rst, mdst_data_rsci_radr_d, mdst_data_rsci_wadr_d, mdst_data_rsci_d_d, mdst_data_rsci_we_d,
      mdst_data_rsci_re_d, mdst_data_rsci_q_d, core_wen, core_wten, mdst_data_rsci_oswt,
      mdst_data_rsci_radr_d_core, mdst_data_rsci_wadr_d_core, mdst_data_rsci_d_d_core,
      mdst_data_rsci_q_d_mxwt, mdst_data_rsci_oswt_pff, mdst_data_rsci_iswt0_1_pff
);
  input clk;
  input rst;
  output [21:0] mdst_data_rsci_radr_d;
  output [21:0] mdst_data_rsci_wadr_d;
  output [19:0] mdst_data_rsci_d_d;
  output mdst_data_rsci_we_d;
  output mdst_data_rsci_re_d;
  input [19:0] mdst_data_rsci_q_d;
  input core_wen;
  input core_wten;
  input mdst_data_rsci_oswt;
  input [21:0] mdst_data_rsci_radr_d_core;
  input [21:0] mdst_data_rsci_wadr_d_core;
  input [19:0] mdst_data_rsci_d_d_core;
  output [19:0] mdst_data_rsci_q_d_mxwt;
  input mdst_data_rsci_oswt_pff;
  input mdst_data_rsci_iswt0_1_pff;


  // Interconnect Declarations
  wire mdst_data_rsci_biwt;
  wire mdst_data_rsci_bdwt;
  wire [21:0] mdst_data_rsci_radr_d_reg;
  wire mdst_data_rsci_radr_d_core_sct_iff;
  wire [21:0] mdst_data_rsci_wadr_d_reg;
  wire mdst_data_rsci_wadr_d_core_sct_iff;
  wire [19:0] mdst_data_rsci_d_d_reg;


  // Interconnect Declarations for Component Instantiations 
  DCT_core_mdst_data_rsci_1_mdst_data_rsc_wait_ctrl DCT_core_mdst_data_rsci_1_mdst_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .mdst_data_rsci_oswt(mdst_data_rsci_oswt),
      .mdst_data_rsci_biwt(mdst_data_rsci_biwt),
      .mdst_data_rsci_bdwt(mdst_data_rsci_bdwt),
      .mdst_data_rsci_radr_d_core_sct_pff(mdst_data_rsci_radr_d_core_sct_iff),
      .mdst_data_rsci_oswt_pff(mdst_data_rsci_oswt_pff),
      .mdst_data_rsci_wadr_d_core_sct_pff(mdst_data_rsci_wadr_d_core_sct_iff),
      .mdst_data_rsci_iswt0_1_pff(mdst_data_rsci_iswt0_1_pff)
    );
  DCT_core_mdst_data_rsci_1_mdst_data_rsc_wait_dp DCT_core_mdst_data_rsci_1_mdst_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .mdst_data_rsci_radr_d(mdst_data_rsci_radr_d_reg),
      .mdst_data_rsci_wadr_d(mdst_data_rsci_wadr_d_reg),
      .mdst_data_rsci_d_d(mdst_data_rsci_d_d_reg),
      .mdst_data_rsci_q_d(mdst_data_rsci_q_d),
      .mdst_data_rsci_radr_d_core(mdst_data_rsci_radr_d_core),
      .mdst_data_rsci_wadr_d_core(mdst_data_rsci_wadr_d_core),
      .mdst_data_rsci_d_d_core(mdst_data_rsci_d_d_core),
      .mdst_data_rsci_q_d_mxwt(mdst_data_rsci_q_d_mxwt),
      .mdst_data_rsci_biwt(mdst_data_rsci_biwt),
      .mdst_data_rsci_bdwt(mdst_data_rsci_bdwt),
      .mdst_data_rsci_radr_d_core_sct(mdst_data_rsci_radr_d_core_sct_iff),
      .mdst_data_rsci_wadr_d_core_sct_pff(mdst_data_rsci_wadr_d_core_sct_iff)
    );
  assign mdst_data_rsci_radr_d = mdst_data_rsci_radr_d_reg;
  assign mdst_data_rsci_wadr_d = mdst_data_rsci_wadr_d_reg;
  assign mdst_data_rsci_d_d = mdst_data_rsci_d_d_reg;
  assign mdst_data_rsci_we_d = mdst_data_rsci_wadr_d_core_sct_iff;
  assign mdst_data_rsci_re_d = mdst_data_rsci_radr_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_src_rsci
// ------------------------------------------------------------------


module DCT_core_src_rsci (
  clk, rst, src_rsc_dat, src_rsc_vld, src_rsc_rdy, core_wen, src_rsci_oswt, src_rsci_wen_comp,
      src_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [19:0] src_rsc_dat;
  input src_rsc_vld;
  output src_rsc_rdy;
  input core_wen;
  input src_rsci_oswt;
  output src_rsci_wen_comp;
  output [19:0] src_rsci_idat_mxwt;


  // Interconnect Declarations
  wire src_rsci_biwt;
  wire src_rsci_bdwt;
  wire src_rsci_bcwt;
  wire src_rsci_irdy_core_sct;
  wire src_rsci_ivld;
  wire [19:0] src_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd2),
  .width(32'sd20)) src_rsci (
      .rdy(src_rsc_rdy),
      .vld(src_rsc_vld),
      .dat(src_rsc_dat),
      .irdy(src_rsci_irdy_core_sct),
      .ivld(src_rsci_ivld),
      .idat(src_rsci_idat)
    );
  DCT_core_src_rsci_src_wait_ctrl DCT_core_src_rsci_src_wait_ctrl_inst (
      .core_wen(core_wen),
      .src_rsci_oswt(src_rsci_oswt),
      .src_rsci_biwt(src_rsci_biwt),
      .src_rsci_bdwt(src_rsci_bdwt),
      .src_rsci_bcwt(src_rsci_bcwt),
      .src_rsci_irdy_core_sct(src_rsci_irdy_core_sct),
      .src_rsci_ivld(src_rsci_ivld)
    );
  DCT_core_src_rsci_src_wait_dp DCT_core_src_rsci_src_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .src_rsci_oswt(src_rsci_oswt),
      .src_rsci_wen_comp(src_rsci_wen_comp),
      .src_rsci_idat_mxwt(src_rsci_idat_mxwt),
      .src_rsci_biwt(src_rsci_biwt),
      .src_rsci_bdwt(src_rsci_bdwt),
      .src_rsci_bcwt(src_rsci_bcwt),
      .src_rsci_idat(src_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core_dst_rsci
// ------------------------------------------------------------------


module DCT_core_dst_rsci (
  clk, rst, dst_rsc_dat, dst_rsc_vld, dst_rsc_rdy, core_wen, dst_rsci_oswt, dst_rsci_wen_comp,
      dst_rsci_idat
);
  input clk;
  input rst;
  output [19:0] dst_rsc_dat;
  output dst_rsc_vld;
  input dst_rsc_rdy;
  input core_wen;
  input dst_rsci_oswt;
  output dst_rsci_wen_comp;
  input [19:0] dst_rsci_idat;


  // Interconnect Declarations
  wire dst_rsci_irdy;
  wire dst_rsci_biwt;
  wire dst_rsci_bdwt;
  wire dst_rsci_bcwt;
  wire dst_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd1),
  .width(32'sd20)) dst_rsci (
      .irdy(dst_rsci_irdy),
      .ivld(dst_rsci_ivld_core_sct),
      .idat(dst_rsci_idat),
      .rdy(dst_rsc_rdy),
      .vld(dst_rsc_vld),
      .dat(dst_rsc_dat)
    );
  DCT_core_dst_rsci_dst_wait_ctrl DCT_core_dst_rsci_dst_wait_ctrl_inst (
      .core_wen(core_wen),
      .dst_rsci_oswt(dst_rsci_oswt),
      .dst_rsci_irdy(dst_rsci_irdy),
      .dst_rsci_biwt(dst_rsci_biwt),
      .dst_rsci_bdwt(dst_rsci_bdwt),
      .dst_rsci_bcwt(dst_rsci_bcwt),
      .dst_rsci_ivld_core_sct(dst_rsci_ivld_core_sct)
    );
  DCT_core_dst_rsci_dst_wait_dp DCT_core_dst_rsci_dst_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dst_rsci_oswt(dst_rsci_oswt),
      .dst_rsci_wen_comp(dst_rsci_wen_comp),
      .dst_rsci_biwt(dst_rsci_biwt),
      .dst_rsci_bdwt(dst_rsci_bdwt),
      .dst_rsci_bcwt(dst_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT_core
// ------------------------------------------------------------------


module DCT_core (
  clk, rst, dst_rsc_dat, dst_rsc_vld, dst_rsc_rdy, src_rsc_dat, src_rsc_vld, src_rsc_rdy,
      mdst_data_rsci_radr_d, mdst_data_rsci_wadr_d, mdst_data_rsci_d_d, mdst_data_rsci_we_d,
      mdst_data_rsci_re_d, mdst_data_rsci_q_d, msrc_data_rsci_radr_d, msrc_data_rsci_wadr_d,
      msrc_data_rsci_d_d, msrc_data_rsci_we_d, msrc_data_rsci_re_d, msrc_data_rsci_q_d
);
  input clk;
  input rst;
  output [19:0] dst_rsc_dat;
  output dst_rsc_vld;
  input dst_rsc_rdy;
  input [19:0] src_rsc_dat;
  input src_rsc_vld;
  output src_rsc_rdy;
  output [21:0] mdst_data_rsci_radr_d;
  output [21:0] mdst_data_rsci_wadr_d;
  output [19:0] mdst_data_rsci_d_d;
  output mdst_data_rsci_we_d;
  output mdst_data_rsci_re_d;
  input [19:0] mdst_data_rsci_q_d;
  output [21:0] msrc_data_rsci_radr_d;
  output [21:0] msrc_data_rsci_wadr_d;
  output [19:0] msrc_data_rsci_d_d;
  output msrc_data_rsci_we_d;
  output msrc_data_rsci_re_d;
  input [19:0] msrc_data_rsci_q_d;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire dst_rsci_wen_comp;
  reg [19:0] dst_rsci_idat;
  wire src_rsci_wen_comp;
  wire [19:0] src_rsci_idat_mxwt;
  wire [19:0] mdst_data_rsci_q_d_mxwt;
  wire [19:0] msrc_data_rsci_q_d_mxwt;
  wire [27:0] fsm_output;
  wire and_dcpl_9;
  wire or_dcpl_38;
  wire and_dcpl_15;
  wire or_dcpl_44;
  wire or_dcpl_55;
  wire or_dcpl_56;
  wire or_tmp_27;
  wire or_tmp_29;
  wire or_tmp_38;
  wire or_tmp_41;
  wire or_tmp_78;
  wire or_tmp_79;
  wire and_141_cse;
  reg [22:0] loop_lmm_i_22_0_sva_1;
  reg [2:0] loop_11_x_3_0_sva_2_0;
  reg loop_11_and_stg_1_1_sva;
  reg loop_11_and_stg_1_2_sva;
  reg loop_11_and_stg_1_3_sva;
  reg loop_11_and_stg_1_0_sva;
  reg [3:0] loop_12_y_3_0_sva_1;
  reg loop_10_m_0_sva;
  reg [2:0] loop_12_y_3_0_sva_2_0;
  reg reg_dst_rsci_oswt_cse;
  reg reg_src_rsci_oswt_cse;
  reg reg_mdst_data_rsci_oswt_cse;
  reg reg_msrc_data_rsci_oswt_cse;
  wire mdst_data_equal_cse;
  wire mdst_data_equal_1_cse;
  wire mdst_data_equal_2_cse;
  wire mdst_data_equal_3_cse;
  wire mdst_data_equal_4_cse;
  wire mdst_data_equal_5_cse;
  wire mdst_data_equal_6_cse;
  wire mdst_data_nor_2_cse;
  wire [21:0] mdst_data_rsci_radr_d_reg;
  wire or_95_rmff;
  wire [21:0] mdst_data_rsci_wadr_d_reg;
  wire [19:0] mdst_data_rsci_d_d_reg;
  wire mdst_data_rsci_we_d_reg;
  wire mdst_data_rsci_re_d_reg;
  wire [21:0] msrc_data_rsci_radr_d_reg;
  wire [21:0] msrc_data_rsci_wadr_d_reg;
  wire [19:0] msrc_data_rsci_d_d_reg;
  wire msrc_data_rsci_we_d_reg;
  wire msrc_data_rsci_re_d_reg;
  reg [7:0] loop_1_i_11_3_sva_7_0;
  reg [7:0] loop_2_j_11_3_sva_7_0;
  reg [1:0] loop_3_k_3_1_sva_1_0;
  reg [19:0] buf_0_lpi_10;
  reg [19:0] buf_1_lpi_10;
  reg [19:0] buf_2_lpi_10;
  reg [19:0] buf_3_lpi_10;
  reg [19:0] buf_4_lpi_10;
  reg [19:0] buf_5_lpi_10;
  reg [19:0] buf_6_lpi_10;
  reg [19:0] buf_7_lpi_10;
  wire or_tmp_101;
  wire [31:0] z_out;
  wire signed [33:0] nl_z_out;
  wire [3:0] z_out_1;
  wire [4:0] nl_z_out_1;
  wire or_tmp_106;
  wire [22:0] z_out_2;
  wire [23:0] nl_z_out_2;
  wire [3:0] z_out_3;
  wire [4:0] nl_z_out_3;
  reg [19:0] loop_12_asn_24_itm;
  reg [13:0] loop_12_mux_9_itm;
  reg loop_12_slc_loop_12_acc_12_3_itm;
  wire loop_lmm_i_22_0_sva_1_mx0c0;
  wire loop_lmm_i_22_0_sva_1_mx0c1;
  wire loop_lmm_i_22_0_sva_1_mx0c2;
  wire loop_3_k_3_1_sva_1_0_mx0c1;
  wire loop_11_x_3_0_sva_2_0_mx0c1;
  wire loop_11_x_3_0_sva_2_0_mx0c2;
  wire loop_11_and_stg_1_3_sva_1;
  wire loop_11_and_stg_1_2_sva_1;
  wire loop_11_and_stg_1_1_sva_1;
  wire loop_1_i_or_cse;
  wire loop_11_and_3_cse;
  wire or_tmp;
  wire or_tmp_111;
  wire mux_tmp;
  wire or_tmp_113;
  wire mux_tmp_2;
  wire or_tmp_115;
  wire mux_tmp_4;
  wire or_tmp_117;
  wire mux_tmp_6;
  wire or_221_tmp;
  wire and_222_tmp;
  wire or_215_tmp;
  wire and_187_tmp;
  wire or_214_tmp;
  wire and_180_tmp;
  wire or_213_tmp;
  wire and_173_tmp;
  wire or_212_tmp;
  wire and_166_tmp;
  wire or_209_tmp;
  wire and_159_tmp;
  wire or_206_tmp;
  wire and_152_tmp;
  wire or_203_tmp;
  wire and_145_tmp;
  wire loop_out_nor_cse;

  wire[0:0] loop_5_loop_5_nand_12_nl;
  wire[0:0] nor_23_nl;
  wire[0:0] loop_5_loop_5_nand_14_nl;
  wire[0:0] nor_24_nl;
  wire[0:0] loop_5_loop_5_nand_16_nl;
  wire[0:0] nor_25_nl;
  wire[0:0] loop_5_loop_5_nand_22_nl;
  wire[0:0] nor_26_nl;
  wire[0:0] loop_5_loop_5_nand_20_nl;
  wire[0:0] nor_27_nl;
  wire[0:0] loop_5_loop_5_nand_18_nl;
  wire[0:0] nor_28_nl;
  wire[0:0] loop_5_loop_5_nand_8_nl;
  wire[0:0] nor_29_nl;
  wire[21:0] loop_lmm_i_loop_lmm_i_and_nl;
  wire[0:0] or_92_nl;
  wire[19:0] loop_6_loop_6_mux1h_nl;
  wire[0:0] loop_6_loop_6_nor_nl;
  wire[0:0] loop_6_and_1_nl;
  wire[0:0] loop_6_and_2_nl;
  wire[0:0] loop_6_and_3_nl;
  wire[0:0] loop_6_and_4_nl;
  wire[0:0] loop_6_and_5_nl;
  wire[0:0] loop_6_and_6_nl;
  wire[0:0] loop_6_and_7_nl;
  wire[0:0] loop_5_loop_5_nand_10_nl;
  wire[0:0] nor_30_nl;
  wire[2:0] loop_11_x_mux1h_3_nl;
  wire[0:0] nor_nl;
  wire[2:0] loop_5_x_mux_1_nl;
  wire[0:0] nand_7_nl;
  wire[13:0] loop_6_mux_9_nl;
  wire[0:0] nor_22_nl;
  wire[0:0] nor_21_nl;
  wire[0:0] nor_20_nl;
  wire[0:0] nor_19_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] mux_16_nl;
  wire[10:0] loop_6_and_9_nl;
  wire[10:0] loop_6_mux1h_6_nl;
  wire[0:0] not_156_nl;
  wire[0:0] loop_6_or_5_nl;
  wire[0:0] loop_6_loop_6_mux_1_nl;
  wire[1:0] loop_6_mux1h_7_nl;
  wire[16:0] loop_6_and_10_nl;
  wire[16:0] loop_6_mux1h_8_nl;
  wire[0:0] not_157_nl;
  wire[0:0] loop_6_mux1h_9_nl;
  wire[1:0] loop_6_mux1h_10_nl;
  wire[0:0] loop_6_mux_12_nl;
  wire[1:0] loop_out_loop_out_and_3_nl;
  wire[1:0] loop_out_mux_2_nl;
  wire[0:0] loop_out_loop_out_and_4_nl;
  wire[10:0] loop_out_loop_out_and_5_nl;
  wire[7:0] loop_out_mux1h_2_nl;
  wire[0:0] loop_out_or_2_nl;
  wire[19:0] loop_out_loop_out_mux_1_nl;
  wire[31:0] operator_40_16_true_AC_TRN_AC_WRAP_mul_3_nl;
  wire signed [33:0] nl_operator_40_16_true_AC_TRN_AC_WRAP_mul_3_nl;
  wire[2:0] loop_12_mux_4_nl;
  wire[0:0] or_222_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[7:0] loop_1_i_mux_nl;
  wire[2:0] loop_12_y_mux_nl;
  wire[7:0] loop_2_j_mux_nl;
  wire[1:0] loop_3_k_mux_nl;
  wire[0:0] loop_10_m_mux_nl;
  wire [21:0] nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_radr_d_core;
  assign loop_1_i_mux_nl = MUX_v_8_2_2(loop_1_i_11_3_sva_7_0, (loop_lmm_i_22_0_sva_1[21:14]),
      fsm_output[25]);
  assign loop_12_y_mux_nl = MUX_v_3_2_2(loop_12_y_3_0_sva_2_0, (loop_lmm_i_22_0_sva_1[13:11]),
      fsm_output[25]);
  assign loop_2_j_mux_nl = MUX_v_8_2_2(loop_2_j_11_3_sva_7_0, (loop_lmm_i_22_0_sva_1[10:3]),
      fsm_output[25]);
  assign loop_3_k_mux_nl = MUX_v_2_2_2(loop_3_k_3_1_sva_1_0, (loop_lmm_i_22_0_sva_1[2:1]),
      fsm_output[25]);
  assign loop_10_m_mux_nl = MUX_s_1_2_2(loop_10_m_0_sva, (loop_lmm_i_22_0_sva_1[0]),
      fsm_output[25]);
  assign nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_radr_d_core = {(loop_1_i_mux_nl)
      , (loop_12_y_mux_nl) , (loop_2_j_mux_nl) , (loop_3_k_mux_nl) , (loop_10_m_mux_nl)};
  wire[1:0] loop_3_k_loop_3_k_and_nl;
  wire[1:0] loop_3_k_mux_1_nl;
  wire[0:0] mdst_data_not_2_nl;
  wire[0:0] loop_10_m_loop_10_m_and_nl;
  wire[0:0] loop_10_m_mux_1_nl;
  wire[1:0] loop_4_loop_4_and_nl;
  wire[1:0] loop_4_mux_nl;
  wire[0:0] mdst_data_not_1_nl;
  wire[0:0] loop_4_l_loop_4_l_and_nl;
  wire[0:0] loop_4_l_mux_1_nl;
  wire [21:0] nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_wadr_d_core;
  assign loop_3_k_mux_1_nl = MUX_v_2_2_2(loop_3_k_3_1_sva_1_0, (loop_11_x_3_0_sva_2_0[2:1]),
      fsm_output[20]);
  assign mdst_data_not_2_nl = ~ or_tmp_27;
  assign loop_3_k_loop_3_k_and_nl = MUX_v_2_2_2(2'b00, (loop_3_k_mux_1_nl), (mdst_data_not_2_nl));
  assign loop_10_m_mux_1_nl = MUX_s_1_2_2(loop_10_m_0_sva, (loop_11_x_3_0_sva_2_0[0]),
      fsm_output[20]);
  assign loop_10_m_loop_10_m_and_nl = (loop_10_m_mux_1_nl) & (~ or_tmp_27);
  assign loop_4_mux_nl = MUX_v_2_2_2((loop_11_x_3_0_sva_2_0[2:1]), loop_3_k_3_1_sva_1_0,
      or_dcpl_38);
  assign mdst_data_not_1_nl = ~ or_tmp_29;
  assign loop_4_loop_4_and_nl = MUX_v_2_2_2(2'b00, (loop_4_mux_nl), (mdst_data_not_1_nl));
  assign loop_4_l_mux_1_nl = MUX_s_1_2_2((loop_11_x_3_0_sva_2_0[0]), loop_10_m_0_sva,
      or_dcpl_38);
  assign loop_4_l_loop_4_l_and_nl = (loop_4_l_mux_1_nl) & (~ or_tmp_29);
  assign nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_wadr_d_core = {loop_1_i_11_3_sva_7_0
      , (loop_3_k_loop_3_k_and_nl) , (loop_10_m_loop_10_m_and_nl) , loop_2_j_11_3_sva_7_0
      , (loop_4_loop_4_and_nl) , (loop_4_l_loop_4_l_and_nl)};
  wire[18:0] mdst_data_mdst_data_mux1h_nl;
  wire[0:0] mdst_data_and_nl;
  wire[0:0] mdst_data_and_1_nl;
  wire[0:0] mdst_data_and_2_nl;
  wire[0:0] mdst_data_and_3_nl;
  wire[0:0] mdst_data_and_4_nl;
  wire[0:0] mdst_data_and_5_nl;
  wire[0:0] mdst_data_and_6_nl;
  wire [19:0] nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_d_d_core;
  assign mdst_data_and_nl = mdst_data_equal_cse & or_tmp_38;
  assign mdst_data_and_1_nl = mdst_data_equal_1_cse & or_tmp_38;
  assign mdst_data_and_2_nl = mdst_data_equal_2_cse & or_tmp_38;
  assign mdst_data_and_3_nl = mdst_data_equal_3_cse & or_tmp_38;
  assign mdst_data_and_4_nl = mdst_data_equal_4_cse & or_tmp_38;
  assign mdst_data_and_5_nl = mdst_data_equal_5_cse & or_tmp_38;
  assign mdst_data_and_6_nl = mdst_data_equal_6_cse & or_tmp_38;
  assign mdst_data_mdst_data_mux1h_nl = MUX1HOT_v_19_8_2((z_out[27:9]), (buf_1_lpi_10[19:1]),
      (buf_2_lpi_10[19:1]), (buf_3_lpi_10[19:1]), (buf_4_lpi_10[19:1]), (buf_5_lpi_10[19:1]),
      (buf_6_lpi_10[19:1]), (buf_7_lpi_10[19:1]), {(~ or_tmp_38) , (mdst_data_and_nl)
      , (mdst_data_and_1_nl) , (mdst_data_and_2_nl) , (mdst_data_and_3_nl) , (mdst_data_and_4_nl)
      , (mdst_data_and_5_nl) , (mdst_data_and_6_nl)});
  assign nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_d_d_core = signext_20_19(mdst_data_mdst_data_mux1h_nl);
  wire [0:0] nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_iswt0_1_pff;
  assign nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_iswt0_1_pff = (fsm_output[10])
      | (fsm_output[8]) | or_dcpl_38;
  wire [21:0] nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_radr_d_core;
  assign nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_radr_d_core = {loop_1_i_11_3_sva_7_0
      , loop_3_k_3_1_sva_1_0 , loop_10_m_0_sva , loop_2_j_11_3_sva_7_0 , loop_12_y_3_0_sva_2_0};
  wire [21:0] nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_wadr_d_core;
  assign nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_wadr_d_core = loop_lmm_i_22_0_sva_1[21:0];
  wire [0:0] nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_oswt_pff;
  assign nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_oswt_pff = fsm_output[4];
  wire [0:0] nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_iswt0_1_pff;
  assign nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_iswt0_1_pff = fsm_output[1];
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_lmm_C_1_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_lmm_C_1_tr0 = loop_lmm_i_22_0_sva_1[22];
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_6_C_2_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_6_C_2_tr0 = loop_12_y_3_0_sva_1[3];
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_5_C_1_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_5_C_1_tr0 = z_out_3[3];
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_7_C_1_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_7_C_1_tr0 = and_dcpl_9;
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_7_C_1_tr1;
  assign nl_DCT_core_core_fsm_inst_loop_7_C_1_tr1 = ~ (loop_12_y_3_0_sva_1[3]);
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_3_C_0_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_3_C_0_tr0 = z_out_2[2];
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_12_C_2_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_12_C_2_tr0 = loop_12_y_3_0_sva_1[3];
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_11_C_1_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_11_C_1_tr0 = z_out_3[3];
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_13_C_1_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_13_C_1_tr0 = and_dcpl_9;
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_13_C_1_tr1;
  assign nl_DCT_core_core_fsm_inst_loop_13_C_1_tr1 = ~ (loop_12_y_3_0_sva_1[3]);
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_9_C_0_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_9_C_0_tr0 = z_out_2[2];
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_2_C_0_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_2_C_0_tr0 = z_out_2[8];
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_1_C_0_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_1_C_0_tr0 = z_out_2[8];
  wire [0:0] nl_DCT_core_core_fsm_inst_loop_out_C_2_tr0;
  assign nl_DCT_core_core_fsm_inst_loop_out_C_2_tr0 = loop_lmm_i_22_0_sva_1[22];
  DCT_core_dst_rsci DCT_core_dst_rsci_inst (
      .clk(clk),
      .rst(rst),
      .dst_rsc_dat(dst_rsc_dat),
      .dst_rsc_vld(dst_rsc_vld),
      .dst_rsc_rdy(dst_rsc_rdy),
      .core_wen(core_wen),
      .dst_rsci_oswt(reg_dst_rsci_oswt_cse),
      .dst_rsci_wen_comp(dst_rsci_wen_comp),
      .dst_rsci_idat(dst_rsci_idat)
    );
  DCT_core_src_rsci DCT_core_src_rsci_inst (
      .clk(clk),
      .rst(rst),
      .src_rsc_dat(src_rsc_dat),
      .src_rsc_vld(src_rsc_vld),
      .src_rsc_rdy(src_rsc_rdy),
      .core_wen(core_wen),
      .src_rsci_oswt(reg_src_rsci_oswt_cse),
      .src_rsci_wen_comp(src_rsci_wen_comp),
      .src_rsci_idat_mxwt(src_rsci_idat_mxwt)
    );
  DCT_core_mdst_data_rsci_1 DCT_core_mdst_data_rsci_1_inst (
      .clk(clk),
      .rst(rst),
      .mdst_data_rsci_radr_d(mdst_data_rsci_radr_d_reg),
      .mdst_data_rsci_wadr_d(mdst_data_rsci_wadr_d_reg),
      .mdst_data_rsci_d_d(mdst_data_rsci_d_d_reg),
      .mdst_data_rsci_we_d(mdst_data_rsci_we_d_reg),
      .mdst_data_rsci_re_d(mdst_data_rsci_re_d_reg),
      .mdst_data_rsci_q_d(mdst_data_rsci_q_d),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .mdst_data_rsci_oswt(reg_mdst_data_rsci_oswt_cse),
      .mdst_data_rsci_radr_d_core(nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_radr_d_core[21:0]),
      .mdst_data_rsci_wadr_d_core(nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_wadr_d_core[21:0]),
      .mdst_data_rsci_d_d_core(nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_d_d_core[19:0]),
      .mdst_data_rsci_q_d_mxwt(mdst_data_rsci_q_d_mxwt),
      .mdst_data_rsci_oswt_pff(or_95_rmff),
      .mdst_data_rsci_iswt0_1_pff(nl_DCT_core_mdst_data_rsci_1_inst_mdst_data_rsci_iswt0_1_pff[0:0])
    );
  DCT_core_msrc_data_rsci_1 DCT_core_msrc_data_rsci_1_inst (
      .clk(clk),
      .rst(rst),
      .msrc_data_rsci_radr_d(msrc_data_rsci_radr_d_reg),
      .msrc_data_rsci_wadr_d(msrc_data_rsci_wadr_d_reg),
      .msrc_data_rsci_d_d(msrc_data_rsci_d_d_reg),
      .msrc_data_rsci_we_d(msrc_data_rsci_we_d_reg),
      .msrc_data_rsci_re_d(msrc_data_rsci_re_d_reg),
      .msrc_data_rsci_q_d(msrc_data_rsci_q_d),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .msrc_data_rsci_oswt(reg_msrc_data_rsci_oswt_cse),
      .msrc_data_rsci_radr_d_core(nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_radr_d_core[21:0]),
      .msrc_data_rsci_wadr_d_core(nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_wadr_d_core[21:0]),
      .msrc_data_rsci_d_d_core(src_rsci_idat_mxwt),
      .msrc_data_rsci_q_d_mxwt(msrc_data_rsci_q_d_mxwt),
      .msrc_data_rsci_oswt_pff(nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_oswt_pff[0:0]),
      .msrc_data_rsci_iswt0_1_pff(nl_DCT_core_msrc_data_rsci_1_inst_msrc_data_rsci_iswt0_1_pff[0:0])
    );
  DCT_core_staller DCT_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dst_rsci_wen_comp(dst_rsci_wen_comp),
      .src_rsci_wen_comp(src_rsci_wen_comp)
    );
  DCT_core_core_fsm DCT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output),
      .loop_lmm_C_1_tr0(nl_DCT_core_core_fsm_inst_loop_lmm_C_1_tr0[0:0]),
      .loop_6_C_2_tr0(nl_DCT_core_core_fsm_inst_loop_6_C_2_tr0[0:0]),
      .loop_5_C_1_tr0(nl_DCT_core_core_fsm_inst_loop_5_C_1_tr0[0:0]),
      .loop_7_C_1_tr0(nl_DCT_core_core_fsm_inst_loop_7_C_1_tr0[0:0]),
      .loop_7_C_1_tr1(nl_DCT_core_core_fsm_inst_loop_7_C_1_tr1[0:0]),
      .loop_3_C_0_tr0(nl_DCT_core_core_fsm_inst_loop_3_C_0_tr0[0:0]),
      .loop_12_C_2_tr0(nl_DCT_core_core_fsm_inst_loop_12_C_2_tr0[0:0]),
      .loop_11_C_1_tr0(nl_DCT_core_core_fsm_inst_loop_11_C_1_tr0[0:0]),
      .loop_13_C_1_tr0(nl_DCT_core_core_fsm_inst_loop_13_C_1_tr0[0:0]),
      .loop_13_C_1_tr1(nl_DCT_core_core_fsm_inst_loop_13_C_1_tr1[0:0]),
      .loop_9_C_0_tr0(nl_DCT_core_core_fsm_inst_loop_9_C_0_tr0[0:0]),
      .loop_2_C_0_tr0(nl_DCT_core_core_fsm_inst_loop_2_C_0_tr0[0:0]),
      .loop_1_C_0_tr0(nl_DCT_core_core_fsm_inst_loop_1_C_0_tr0[0:0]),
      .loop_out_C_2_tr0(nl_DCT_core_core_fsm_inst_loop_out_C_2_tr0[0:0])
    );
  assign or_95_rmff = (fsm_output[14]) | (fsm_output[25]);
  assign mdst_data_equal_cse = (loop_11_x_3_0_sva_2_0==3'b001);
  assign mdst_data_equal_1_cse = (loop_11_x_3_0_sva_2_0==3'b010);
  assign mdst_data_equal_2_cse = (loop_11_x_3_0_sva_2_0==3'b011);
  assign mdst_data_nor_2_cse = ~((loop_11_x_3_0_sva_2_0[1:0]!=2'b00));
  assign mdst_data_equal_3_cse = (loop_11_x_3_0_sva_2_0[2]) & mdst_data_nor_2_cse;
  assign mdst_data_equal_4_cse = (loop_11_x_3_0_sva_2_0==3'b101);
  assign mdst_data_equal_5_cse = (loop_11_x_3_0_sva_2_0==3'b110);
  assign mdst_data_equal_6_cse = (loop_11_x_3_0_sva_2_0==3'b111);
  assign loop_1_i_or_cse = (fsm_output[2]) | (fsm_output[24]);
  assign loop_11_and_3_cse = core_wen & (~(or_dcpl_56 | (fsm_output[4]) | (fsm_output[14])
      | (fsm_output[6]) | (fsm_output[16])));
  assign loop_11_and_stg_1_3_sva_1 = (loop_11_x_3_0_sva_2_0[1:0]==2'b11);
  assign loop_11_and_stg_1_2_sva_1 = (loop_11_x_3_0_sva_2_0[1:0]==2'b10);
  assign loop_11_and_stg_1_1_sva_1 = (loop_11_x_3_0_sva_2_0[1:0]==2'b01);
  assign and_dcpl_9 = (loop_12_y_3_0_sva_1[3]) & loop_10_m_0_sva;
  assign or_dcpl_38 = (fsm_output[20]) | (fsm_output[18]);
  assign and_dcpl_15 = ~((fsm_output[6]) | (fsm_output[16]));
  assign or_dcpl_44 = (fsm_output[6]) | (fsm_output[16]);
  assign or_dcpl_55 = (fsm_output[4]) | (fsm_output[14]);
  assign or_dcpl_56 = (fsm_output[5]) | (fsm_output[15]);
  assign or_tmp_27 = ~((fsm_output[10]) | (fsm_output[8]) | (fsm_output[20]));
  assign or_tmp_29 = ~((fsm_output[10]) | (fsm_output[20]) | (fsm_output[18]));
  assign or_tmp_38 = (fsm_output[10]) | (fsm_output[20]);
  assign or_tmp_41 = (fsm_output[13]) | (fsm_output[3]);
  assign and_141_cse = (~((fsm_output[13]) | (fsm_output[3]))) & and_dcpl_15;
  assign or_tmp_78 = (fsm_output[22]) | (fsm_output[12]) | (fsm_output[24]) | (fsm_output[23])
      | (fsm_output[2]);
  assign or_tmp_79 = (fsm_output[11]) | (fsm_output[21]);
  assign loop_lmm_i_22_0_sva_1_mx0c0 = (fsm_output[1]) | (fsm_output[25]);
  assign loop_lmm_i_22_0_sva_1_mx0c1 = (fsm_output[0]) | (fsm_output[27]) | loop_1_i_or_cse;
  assign loop_lmm_i_22_0_sva_1_mx0c2 = or_dcpl_56 | or_dcpl_55;
  assign loop_3_k_3_1_sva_1_0_mx0c1 = (fsm_output[22]) | ((~ (z_out_2[2])) & (fsm_output[12]));
  assign loop_11_x_3_0_sva_2_0_mx0c1 = (fsm_output[7]) | (fsm_output[17]);
  assign loop_11_x_3_0_sva_2_0_mx0c2 = (fsm_output[9]) | (fsm_output[19]);
  assign mdst_data_rsci_radr_d = mdst_data_rsci_radr_d_reg;
  assign mdst_data_rsci_wadr_d = mdst_data_rsci_wadr_d_reg;
  assign mdst_data_rsci_d_d = mdst_data_rsci_d_d_reg;
  assign mdst_data_rsci_we_d = mdst_data_rsci_we_d_reg;
  assign mdst_data_rsci_re_d = mdst_data_rsci_re_d_reg;
  assign msrc_data_rsci_radr_d = msrc_data_rsci_radr_d_reg;
  assign msrc_data_rsci_wadr_d = msrc_data_rsci_wadr_d_reg;
  assign msrc_data_rsci_d_d = msrc_data_rsci_d_d_reg;
  assign msrc_data_rsci_we_d = msrc_data_rsci_we_d_reg;
  assign msrc_data_rsci_re_d = msrc_data_rsci_re_d_reg;
  assign or_tmp_101 = (fsm_output[18]) | (fsm_output[8]);
  assign or_tmp_106 = (fsm_output[22]) | (fsm_output[12]);
  assign or_tmp = or_tmp_41 | or_dcpl_44;
  assign or_tmp_111 = loop_11_and_stg_1_1_sva | (~ or_dcpl_44);
  assign nor_22_nl = ~(or_tmp_41 | (~ or_tmp_111));
  assign mux_tmp = MUX_s_1_2_2((nor_22_nl), or_tmp_111, loop_11_and_stg_1_1_sva_1);
  assign or_tmp_113 = loop_11_and_stg_1_2_sva | (~ or_dcpl_44);
  assign nor_21_nl = ~(or_tmp_41 | (~ or_tmp_113));
  assign mux_tmp_2 = MUX_s_1_2_2((nor_21_nl), or_tmp_113, loop_11_and_stg_1_2_sva_1);
  assign or_tmp_115 = loop_11_and_stg_1_3_sva | (~ or_dcpl_44);
  assign nor_20_nl = ~(or_tmp_41 | (~ or_tmp_115));
  assign mux_tmp_4 = MUX_s_1_2_2((nor_20_nl), or_tmp_115, loop_11_and_stg_1_3_sva_1);
  assign or_tmp_117 = loop_11_and_stg_1_0_sva | (~ or_dcpl_44);
  assign nor_19_nl = ~(or_tmp_41 | (~ or_tmp_117));
  assign mux_tmp_6 = MUX_s_1_2_2((nor_19_nl), or_tmp_117, mdst_data_nor_2_cse);
  assign mux_6_nl = MUX_s_1_2_2((~ mux_tmp), or_tmp, loop_11_x_3_0_sva_2_0[2]);
  assign or_203_tmp = (mux_6_nl) | and_141_cse;
  assign and_145_tmp = loop_11_and_stg_1_1_sva & (~ (loop_11_x_3_0_sva_2_0[2])) &
      or_dcpl_44;
  assign mux_8_nl = MUX_s_1_2_2((~ mux_tmp_2), or_tmp, loop_11_x_3_0_sva_2_0[2]);
  assign or_206_tmp = (mux_8_nl) | and_141_cse;
  assign and_152_tmp = loop_11_and_stg_1_2_sva & (~ (loop_11_x_3_0_sva_2_0[2])) &
      or_dcpl_44;
  assign mux_10_nl = MUX_s_1_2_2((~ mux_tmp_4), or_tmp, loop_11_x_3_0_sva_2_0[2]);
  assign or_209_tmp = (mux_10_nl) | and_141_cse;
  assign and_159_tmp = loop_11_and_stg_1_3_sva & (~ (loop_11_x_3_0_sva_2_0[2])) &
      or_dcpl_44;
  assign mux_12_nl = MUX_s_1_2_2(or_tmp, (~ mux_tmp_6), loop_11_x_3_0_sva_2_0[2]);
  assign or_212_tmp = (mux_12_nl) | and_141_cse;
  assign and_166_tmp = loop_11_and_stg_1_0_sva & (loop_11_x_3_0_sva_2_0[2]) & or_dcpl_44;
  assign mux_13_nl = MUX_s_1_2_2(or_tmp, (~ mux_tmp), loop_11_x_3_0_sva_2_0[2]);
  assign or_213_tmp = (mux_13_nl) | and_141_cse;
  assign and_173_tmp = loop_11_and_stg_1_1_sva & (loop_11_x_3_0_sva_2_0[2]) & or_dcpl_44;
  assign mux_14_nl = MUX_s_1_2_2(or_tmp, (~ mux_tmp_2), loop_11_x_3_0_sva_2_0[2]);
  assign or_214_tmp = (mux_14_nl) | and_141_cse;
  assign and_180_tmp = loop_11_and_stg_1_2_sva & (loop_11_x_3_0_sva_2_0[2]) & or_dcpl_44;
  assign mux_15_nl = MUX_s_1_2_2(or_tmp, (~ mux_tmp_4), loop_11_x_3_0_sva_2_0[2]);
  assign or_215_tmp = (mux_15_nl) | and_141_cse;
  assign and_187_tmp = loop_11_and_stg_1_3_sva & (loop_11_x_3_0_sva_2_0[2]) & or_dcpl_44;
  assign mux_16_nl = MUX_s_1_2_2((~ mux_tmp_6), or_tmp, loop_11_x_3_0_sva_2_0[2]);
  assign or_221_tmp = (mux_16_nl) | or_dcpl_56 | (fsm_output[4]) | (fsm_output[7])
      | (fsm_output[14]) | (fsm_output[17]);
  assign and_222_tmp = loop_11_and_stg_1_0_sva & (~ (loop_11_x_3_0_sva_2_0[2])) &
      or_dcpl_44;
  assign loop_out_nor_cse = ~(or_tmp_106 | (fsm_output[24:23]!=2'b00));
  always @(posedge clk) begin
    if ( core_wen & (fsm_output[26]) ) begin
      dst_rsci_idat <= mdst_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( core_wen ) begin
      buf_1_lpi_10 <= MUX1HOT_v_20_3_2((signext_20_1(loop_5_loop_5_nand_12_nl)),
          (z_out_2[19:0]), buf_1_lpi_10, {(nor_23_nl) , and_145_tmp , or_203_tmp});
      buf_2_lpi_10 <= MUX1HOT_v_20_3_2((signext_20_1(loop_5_loop_5_nand_14_nl)),
          (z_out_2[19:0]), buf_2_lpi_10, {(nor_24_nl) , and_152_tmp , or_206_tmp});
      buf_3_lpi_10 <= MUX1HOT_v_20_3_2((signext_20_1(loop_5_loop_5_nand_16_nl)),
          (z_out_2[19:0]), buf_3_lpi_10, {(nor_25_nl) , and_159_tmp , or_209_tmp});
      buf_4_lpi_10 <= MUX1HOT_v_20_3_2((signext_20_1(loop_5_loop_5_nand_22_nl)),
          (z_out_2[19:0]), buf_4_lpi_10, {(nor_26_nl) , and_166_tmp , or_212_tmp});
      buf_5_lpi_10 <= MUX1HOT_v_20_3_2((signext_20_1(loop_5_loop_5_nand_20_nl)),
          (z_out_2[19:0]), buf_5_lpi_10, {(nor_27_nl) , and_173_tmp , or_213_tmp});
      buf_6_lpi_10 <= MUX1HOT_v_20_3_2((signext_20_1(loop_5_loop_5_nand_18_nl)),
          (z_out_2[19:0]), buf_6_lpi_10, {(nor_28_nl) , and_180_tmp , or_214_tmp});
      buf_7_lpi_10 <= MUX1HOT_v_20_3_2((signext_20_1(loop_5_loop_5_nand_8_nl)), (z_out_2[19:0]),
          buf_7_lpi_10, {(nor_29_nl) , and_187_tmp , or_215_tmp});
      buf_0_lpi_10 <= MUX1HOT_v_20_3_2((signext_20_1(loop_5_loop_5_nand_10_nl)),
          (z_out_2[19:0]), buf_0_lpi_10, {(nor_30_nl) , and_222_tmp , or_221_tmp});
      loop_12_y_3_0_sva_2_0 <= MUX_v_3_2_2(3'b000, (loop_5_x_mux_1_nl), (nand_7_nl));
      loop_12_mux_9_itm <= MUX_v_14_2_2((loop_6_mux_9_nl), loop_12_mux_9_itm, or_dcpl_56);
      loop_12_asn_24_itm <= MUX_v_20_2_2(msrc_data_rsci_q_d_mxwt, mdst_data_rsci_q_d_mxwt,
          fsm_output[15]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_dst_rsci_oswt_cse <= 1'b0;
      reg_src_rsci_oswt_cse <= 1'b0;
      reg_mdst_data_rsci_oswt_cse <= 1'b0;
      reg_msrc_data_rsci_oswt_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_dst_rsci_oswt_cse <= fsm_output[26];
      reg_src_rsci_oswt_cse <= ~((~((fsm_output[0]) | (fsm_output[2]))) | ((loop_lmm_i_22_0_sva_1[22])
          & (fsm_output[2])));
      reg_mdst_data_rsci_oswt_cse <= or_95_rmff;
      reg_msrc_data_rsci_oswt_cse <= fsm_output[4];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      loop_lmm_i_22_0_sva_1 <= 23'b00000000000000000000000;
    end
    else if ( core_wen & (loop_lmm_i_22_0_sva_1_mx0c0 | loop_lmm_i_22_0_sva_1_mx0c1
        | loop_lmm_i_22_0_sva_1_mx0c2) ) begin
      loop_lmm_i_22_0_sva_1 <= MUX1HOT_v_23_3_2(z_out_2, ({1'b0 , (loop_lmm_i_loop_lmm_i_and_nl)}),
          ({3'b000 , (loop_6_loop_6_mux1h_nl)}), {loop_lmm_i_22_0_sva_1_mx0c0 , loop_lmm_i_22_0_sva_1_mx0c1
          , loop_lmm_i_22_0_sva_1_mx0c2});
    end
  end
  always @(posedge clk) begin
    if ( core_wen & loop_1_i_or_cse ) begin
      loop_1_i_11_3_sva_7_0 <= MUX_v_8_2_2(8'b00000000, (z_out_2[7:0]), (fsm_output[24]));
    end
  end
  always @(posedge clk) begin
    if ( core_wen & (loop_1_i_or_cse | (fsm_output[23])) ) begin
      loop_2_j_11_3_sva_7_0 <= MUX_v_8_2_2(8'b00000000, (z_out_2[7:0]), (fsm_output[23]));
    end
  end
  always @(posedge clk) begin
    if ( core_wen & ((fsm_output[24]) | (fsm_output[23]) | (fsm_output[2]) | ((z_out_2[2])
        & (fsm_output[12])) | loop_3_k_3_1_sva_1_0_mx0c1) ) begin
      loop_3_k_3_1_sva_1_0 <= MUX_v_2_2_2(2'b00, (z_out_2[1:0]), loop_3_k_3_1_sva_1_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      loop_10_m_0_sva <= 1'b0;
    end
    else if ( core_wen & (or_tmp_78 | or_tmp_79) ) begin
      loop_10_m_0_sva <= (loop_10_m_0_sva | (loop_12_y_3_0_sva_1[3])) & or_tmp_79;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      loop_11_x_3_0_sva_2_0 <= 3'b000;
    end
    else if ( core_wen & (or_tmp_78 | loop_11_x_3_0_sva_2_0_mx0c1 | loop_11_x_3_0_sva_2_0_mx0c2
        | or_tmp_79) ) begin
      loop_11_x_3_0_sva_2_0 <= MUX_v_3_2_2(3'b000, (loop_11_x_mux1h_3_nl), (nor_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      loop_11_and_stg_1_0_sva <= 1'b0;
      loop_11_and_stg_1_1_sva <= 1'b0;
      loop_11_and_stg_1_2_sva <= 1'b0;
      loop_11_and_stg_1_3_sva <= 1'b0;
    end
    else if ( loop_11_and_3_cse ) begin
      loop_11_and_stg_1_0_sva <= mdst_data_nor_2_cse;
      loop_11_and_stg_1_1_sva <= loop_11_and_stg_1_1_sva_1;
      loop_11_and_stg_1_2_sva <= loop_11_and_stg_1_2_sva_1;
      loop_11_and_stg_1_3_sva <= loop_11_and_stg_1_3_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      loop_12_y_3_0_sva_1 <= 4'b0000;
    end
    else if ( core_wen & (or_dcpl_55 | or_tmp_38) ) begin
      loop_12_y_3_0_sva_1 <= z_out_3;
    end
  end
  always @(posedge clk) begin
    if ( core_wen & (loop_11_and_stg_1_3_sva | loop_11_and_stg_1_0_sva | loop_11_and_stg_1_2_sva
        | loop_11_and_stg_1_1_sva) ) begin
      loop_12_slc_loop_12_acc_12_3_itm <= z_out_1[3];
    end
  end
  assign loop_5_loop_5_nand_12_nl = ~(loop_11_and_stg_1_1_sva_1 & (~ (loop_11_x_3_0_sva_2_0[2])));
  assign nor_23_nl = ~(and_145_tmp | or_203_tmp);
  assign loop_5_loop_5_nand_14_nl = ~(loop_11_and_stg_1_2_sva_1 & (~ (loop_11_x_3_0_sva_2_0[2])));
  assign nor_24_nl = ~(and_152_tmp | or_206_tmp);
  assign loop_5_loop_5_nand_16_nl = ~(loop_11_and_stg_1_3_sva_1 & (~ (loop_11_x_3_0_sva_2_0[2])));
  assign nor_25_nl = ~(and_159_tmp | or_209_tmp);
  assign loop_5_loop_5_nand_22_nl = ~(mdst_data_nor_2_cse & (loop_11_x_3_0_sva_2_0[2]));
  assign nor_26_nl = ~(and_166_tmp | or_212_tmp);
  assign loop_5_loop_5_nand_20_nl = ~(loop_11_and_stg_1_1_sva_1 & (loop_11_x_3_0_sva_2_0[2]));
  assign nor_27_nl = ~(and_173_tmp | or_213_tmp);
  assign loop_5_loop_5_nand_18_nl = ~(loop_11_and_stg_1_2_sva_1 & (loop_11_x_3_0_sva_2_0[2]));
  assign nor_28_nl = ~(and_180_tmp | or_214_tmp);
  assign loop_5_loop_5_nand_8_nl = ~(loop_11_and_stg_1_3_sva_1 & (loop_11_x_3_0_sva_2_0[2]));
  assign nor_29_nl = ~(and_187_tmp | or_215_tmp);
  assign loop_5_loop_5_nand_10_nl = ~(mdst_data_nor_2_cse & (~ (loop_11_x_3_0_sva_2_0[2])));
  assign nor_30_nl = ~(and_222_tmp | or_221_tmp);
  assign loop_5_x_mux_1_nl = MUX_v_3_2_2(loop_12_y_3_0_sva_2_0, (loop_12_y_3_0_sva_1[2:0]),
      or_dcpl_44);
  assign nand_7_nl = ~((~((fsm_output[4]) | (fsm_output[14]))) & and_dcpl_15);
  assign loop_6_mux_9_nl = MUX_v_14_16_2(14'b01000000000000, 14'b00111110110001,
      14'b00111011001000, 14'b00110101001101, 14'b00101101010000, 14'b00100011100011,
      14'b00011000011111, 14'b00001100011111, 14'b00000000000000, 14'b11110011100000,
      14'b11100111100000, 14'b11011100011100, 14'b11010010101111, 14'b11001010110010,
      14'b11000100110111, 14'b11000001001110, {(z_out_1[2:0]) , (loop_11_x_3_0_sva_2_0[0])});
  assign or_92_nl = (fsm_output[27]) | (fsm_output[2]);
  assign loop_lmm_i_loop_lmm_i_and_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      (loop_lmm_i_22_0_sva_1[21:0]), (or_92_nl));
  assign loop_6_loop_6_nor_nl = ~((loop_11_x_3_0_sva_2_0!=3'b000) | or_dcpl_56);
  assign loop_6_and_1_nl = mdst_data_equal_cse & (~ or_dcpl_56);
  assign loop_6_and_2_nl = mdst_data_equal_1_cse & (~ or_dcpl_56);
  assign loop_6_and_3_nl = mdst_data_equal_2_cse & (~ or_dcpl_56);
  assign loop_6_and_4_nl = mdst_data_equal_3_cse & (~ or_dcpl_56);
  assign loop_6_and_5_nl = mdst_data_equal_4_cse & (~ or_dcpl_56);
  assign loop_6_and_6_nl = mdst_data_equal_5_cse & (~ or_dcpl_56);
  assign loop_6_and_7_nl = mdst_data_equal_6_cse & (~ or_dcpl_56);
  assign loop_6_loop_6_mux1h_nl = MUX1HOT_v_20_9_2(buf_0_lpi_10, buf_1_lpi_10, buf_2_lpi_10,
      buf_3_lpi_10, buf_4_lpi_10, buf_5_lpi_10, buf_6_lpi_10, buf_7_lpi_10, (loop_lmm_i_22_0_sva_1[19:0]),
      {(loop_6_loop_6_nor_nl) , (loop_6_and_1_nl) , (loop_6_and_2_nl) , (loop_6_and_3_nl)
      , (loop_6_and_4_nl) , (loop_6_and_5_nl) , (loop_6_and_6_nl) , (loop_6_and_7_nl)
      , or_dcpl_56});
  assign loop_11_x_mux1h_3_nl = MUX1HOT_v_3_3_2((z_out_3[2:0]), 3'b001, (loop_12_y_3_0_sva_1[2:0]),
      {loop_11_x_3_0_sva_2_0_mx0c1 , loop_11_x_3_0_sva_2_0_mx0c2 , or_tmp_79});
  assign nor_nl = ~((or_tmp_79 & (loop_12_y_3_0_sva_1[3])) | or_tmp_78);
  assign loop_6_mux1h_6_nl = MUX1HOT_v_11_3_2((signext_11_1(loop_12_y_3_0_sva_2_0[2])),
      (loop_12_mux_9_itm[13:3]), 11'b00000010110, {or_dcpl_55 , or_dcpl_44 , or_tmp_101});
  assign not_156_nl = ~ or_dcpl_56;
  assign loop_6_and_9_nl = MUX_v_11_2_2(11'b00000000000, (loop_6_mux1h_6_nl), (not_156_nl));
  assign loop_6_loop_6_mux_1_nl = MUX_s_1_2_2((loop_12_y_3_0_sva_2_0[2]), (loop_12_mux_9_itm[2]),
      or_dcpl_44);
  assign loop_6_or_5_nl = (loop_6_loop_6_mux_1_nl) | or_tmp_101;
  assign loop_6_mux1h_7_nl = MUX1HOT_v_2_3_2((loop_12_y_3_0_sva_2_0[1:0]), (loop_12_mux_9_itm[1:0]),
      2'b01, {loop_lmm_i_22_0_sva_1_mx0c2 , or_dcpl_44 , or_tmp_101});
  assign loop_6_mux1h_8_nl = MUX1HOT_v_17_3_2((signext_17_1(loop_11_x_3_0_sva_2_0[2])),
      (loop_12_asn_24_itm[19:3]), (buf_0_lpi_10[19:3]), {or_dcpl_55 , or_dcpl_44
      , or_tmp_101});
  assign not_157_nl = ~ or_dcpl_56;
  assign loop_6_and_10_nl = MUX_v_17_2_2(17'b00000000000000000, (loop_6_mux1h_8_nl),
      (not_157_nl));
  assign loop_6_mux1h_9_nl = MUX1HOT_s_1_3_2((loop_11_x_3_0_sva_2_0[2]), (loop_12_asn_24_itm[2]),
      (buf_0_lpi_10[2]), {loop_lmm_i_22_0_sva_1_mx0c2 , or_dcpl_44 , or_tmp_101});
  assign loop_6_mux1h_10_nl = MUX1HOT_v_2_3_2((loop_11_x_3_0_sva_2_0[1:0]), (loop_12_asn_24_itm[1:0]),
      (buf_0_lpi_10[1:0]), {loop_lmm_i_22_0_sva_1_mx0c2 , or_dcpl_44 , or_tmp_101});
  assign nl_z_out = $signed(({(loop_6_and_9_nl) , (loop_6_or_5_nl) , (loop_6_mux1h_7_nl)}))
      * $signed(({(loop_6_and_10_nl) , (loop_6_mux1h_9_nl) , (loop_6_mux1h_10_nl)}));
  assign z_out = nl_z_out[31:0];
  assign loop_6_mux_12_nl = MUX_s_1_2_2((z_out[2]), (z_out[3]), or_dcpl_56);
  assign nl_z_out_1 = ({(loop_6_mux_12_nl) , (z_out[2:0])}) + conv_u2u_2_4(loop_11_x_3_0_sva_2_0[2:1]);
  assign z_out_1 = nl_z_out_1[3:0];
  assign loop_out_mux_2_nl = MUX_v_2_2_2((loop_lmm_i_22_0_sva_1[21:20]), (signext_2_1(loop_lmm_i_22_0_sva_1[19])),
      or_dcpl_44);
  assign loop_out_loop_out_and_3_nl = MUX_v_2_2_2(2'b00, (loop_out_mux_2_nl), loop_out_nor_cse);
  assign loop_out_loop_out_and_4_nl = (loop_lmm_i_22_0_sva_1[19]) & loop_out_nor_cse;
  assign loop_out_loop_out_and_5_nl = MUX_v_11_2_2(11'b00000000000, (loop_lmm_i_22_0_sva_1[18:8]),
      loop_out_nor_cse);
  assign loop_out_or_2_nl = loop_lmm_i_22_0_sva_1_mx0c0 | or_dcpl_44;
  assign loop_out_mux1h_2_nl = MUX1HOT_v_8_4_2((loop_lmm_i_22_0_sva_1[7:0]), ({6'b000000
      , loop_3_k_3_1_sva_1_0}), loop_2_j_11_3_sva_7_0, loop_1_i_11_3_sva_7_0, {(loop_out_or_2_nl)
      , or_tmp_106 , (fsm_output[23]) , (fsm_output[24])});
  assign nl_operator_40_16_true_AC_TRN_AC_WRAP_mul_3_nl = $signed(z_out) * $signed(({loop_12_slc_loop_12_acc_12_3_itm
      , 1'b1}));
  assign operator_40_16_true_AC_TRN_AC_WRAP_mul_3_nl = nl_operator_40_16_true_AC_TRN_AC_WRAP_mul_3_nl[31:0];
  assign loop_out_loop_out_mux_1_nl = MUX_v_20_2_2(20'b00000000000000000001, (readslicef_32_20_12((operator_40_16_true_AC_TRN_AC_WRAP_mul_3_nl))),
      or_dcpl_44);
  assign nl_z_out_2 = conv_u2u_22_23({(loop_out_loop_out_and_3_nl) , (loop_out_loop_out_and_4_nl)
      , (loop_out_loop_out_and_5_nl) , (loop_out_mux1h_2_nl)}) + conv_u2u_20_23(loop_out_loop_out_mux_1_nl);
  assign z_out_2 = nl_z_out_2[22:0];
  assign or_222_nl = (fsm_output[20]) | (fsm_output[17]) | (fsm_output[10]) | (fsm_output[7]);
  assign loop_12_mux_4_nl = MUX_v_3_2_2(loop_12_y_3_0_sva_2_0, loop_11_x_3_0_sva_2_0,
      or_222_nl);
  assign nl_z_out_3 = conv_u2u_3_4(loop_12_mux_4_nl) + 4'b0001;
  assign z_out_3 = nl_z_out_3[3:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction


  function automatic [16:0] MUX1HOT_v_17_3_2;
    input [16:0] input_2;
    input [16:0] input_1;
    input [16:0] input_0;
    input [2:0] sel;
    reg [16:0] result;
  begin
    result = input_0 & {17{sel[0]}};
    result = result | ( input_1 & {17{sel[1]}});
    result = result | ( input_2 & {17{sel[2]}});
    MUX1HOT_v_17_3_2 = result;
  end
  endfunction


  function automatic [18:0] MUX1HOT_v_19_8_2;
    input [18:0] input_7;
    input [18:0] input_6;
    input [18:0] input_5;
    input [18:0] input_4;
    input [18:0] input_3;
    input [18:0] input_2;
    input [18:0] input_1;
    input [18:0] input_0;
    input [7:0] sel;
    reg [18:0] result;
  begin
    result = input_0 & {19{sel[0]}};
    result = result | ( input_1 & {19{sel[1]}});
    result = result | ( input_2 & {19{sel[2]}});
    result = result | ( input_3 & {19{sel[3]}});
    result = result | ( input_4 & {19{sel[4]}});
    result = result | ( input_5 & {19{sel[5]}});
    result = result | ( input_6 & {19{sel[6]}});
    result = result | ( input_7 & {19{sel[7]}});
    MUX1HOT_v_19_8_2 = result;
  end
  endfunction


  function automatic [19:0] MUX1HOT_v_20_3_2;
    input [19:0] input_2;
    input [19:0] input_1;
    input [19:0] input_0;
    input [2:0] sel;
    reg [19:0] result;
  begin
    result = input_0 & {20{sel[0]}};
    result = result | ( input_1 & {20{sel[1]}});
    result = result | ( input_2 & {20{sel[2]}});
    MUX1HOT_v_20_3_2 = result;
  end
  endfunction


  function automatic [19:0] MUX1HOT_v_20_9_2;
    input [19:0] input_8;
    input [19:0] input_7;
    input [19:0] input_6;
    input [19:0] input_5;
    input [19:0] input_4;
    input [19:0] input_3;
    input [19:0] input_2;
    input [19:0] input_1;
    input [19:0] input_0;
    input [8:0] sel;
    reg [19:0] result;
  begin
    result = input_0 & {20{sel[0]}};
    result = result | ( input_1 & {20{sel[1]}});
    result = result | ( input_2 & {20{sel[2]}});
    result = result | ( input_3 & {20{sel[3]}});
    result = result | ( input_4 & {20{sel[4]}});
    result = result | ( input_5 & {20{sel[5]}});
    result = result | ( input_6 & {20{sel[6]}});
    result = result | ( input_7 & {20{sel[7]}});
    result = result | ( input_8 & {20{sel[8]}});
    MUX1HOT_v_20_9_2 = result;
  end
  endfunction


  function automatic [22:0] MUX1HOT_v_23_3_2;
    input [22:0] input_2;
    input [22:0] input_1;
    input [22:0] input_0;
    input [2:0] sel;
    reg [22:0] result;
  begin
    result = input_0 & {23{sel[0]}};
    result = result | ( input_1 & {23{sel[1]}});
    result = result | ( input_2 & {23{sel[2]}});
    MUX1HOT_v_23_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_16_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [13:0] input_2;
    input [13:0] input_3;
    input [13:0] input_4;
    input [13:0] input_5;
    input [13:0] input_6;
    input [13:0] input_7;
    input [13:0] input_8;
    input [13:0] input_9;
    input [13:0] input_10;
    input [13:0] input_11;
    input [13:0] input_12;
    input [13:0] input_13;
    input [13:0] input_14;
    input [13:0] input_15;
    input [3:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_14_16_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [0:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [19:0] readslicef_32_20_12;
    input [31:0] vector;
    reg [31:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_32_20_12 = tmp[19:0];
  end
  endfunction


  function automatic [10:0] signext_11_1;
    input [0:0] vector;
  begin
    signext_11_1= {{10{vector[0]}}, vector};
  end
  endfunction


  function automatic [16:0] signext_17_1;
    input [0:0] vector;
  begin
    signext_17_1= {{16{vector[0]}}, vector};
  end
  endfunction


  function automatic [19:0] signext_20_1;
    input [0:0] vector;
  begin
    signext_20_1= {{19{vector[0]}}, vector};
  end
  endfunction


  function automatic [19:0] signext_20_19;
    input [18:0] vector;
  begin
    signext_20_19= {{1{vector[18]}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [22:0] conv_u2u_20_23 ;
    input [19:0]  vector ;
  begin
    conv_u2u_20_23 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [22:0] conv_u2u_22_23 ;
    input [21:0]  vector ;
  begin
    conv_u2u_22_23 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    DCT
// ------------------------------------------------------------------


module DCT (
  clk, rst, dst_rsc_dat, dst_rsc_vld, dst_rsc_rdy, src_rsc_dat, src_rsc_vld, src_rsc_rdy
);
  input clk;
  input rst;
  output [19:0] dst_rsc_dat;
  output dst_rsc_vld;
  input dst_rsc_rdy;
  input [19:0] src_rsc_dat;
  input src_rsc_vld;
  output src_rsc_rdy;


  // Interconnect Declarations
  wire [21:0] mdst_data_rsci_radr_d;
  wire [21:0] mdst_data_rsci_wadr_d;
  wire [19:0] mdst_data_rsci_d_d;
  wire mdst_data_rsci_we_d;
  wire mdst_data_rsci_re_d;
  wire [19:0] mdst_data_rsci_q_d;
  wire [21:0] msrc_data_rsci_radr_d;
  wire [21:0] msrc_data_rsci_wadr_d;
  wire [19:0] msrc_data_rsci_d_d;
  wire msrc_data_rsci_we_d;
  wire msrc_data_rsci_re_d;
  wire [19:0] msrc_data_rsci_q_d;
  wire mdst_data_rsc_we;
  wire [19:0] mdst_data_rsc_d;
  wire [21:0] mdst_data_rsc_wadr;
  wire mdst_data_rsc_re;
  wire [19:0] mdst_data_rsc_q;
  wire [21:0] mdst_data_rsc_radr;
  wire msrc_data_rsc_we;
  wire [19:0] msrc_data_rsc_d;
  wire [21:0] msrc_data_rsc_wadr;
  wire msrc_data_rsc_re;
  wire [19:0] msrc_data_rsc_q;
  wire [21:0] msrc_data_rsc_radr;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.data_width(32'sd20),
  .addr_width(32'sd22),
  .depth(32'sd4194304)) mdst_data_rsc_comp (
      .radr(mdst_data_rsc_radr),
      .wadr(mdst_data_rsc_wadr),
      .d(mdst_data_rsc_d),
      .we(mdst_data_rsc_we),
      .re(mdst_data_rsc_re),
      .clk(clk),
      .q(mdst_data_rsc_q)
    );
  BLOCK_1R1W_RBW #(.data_width(32'sd20),
  .addr_width(32'sd22),
  .depth(32'sd4194304)) msrc_data_rsc_comp (
      .radr(msrc_data_rsc_radr),
      .wadr(msrc_data_rsc_wadr),
      .d(msrc_data_rsc_d),
      .we(msrc_data_rsc_we),
      .re(msrc_data_rsc_re),
      .clk(clk),
      .q(msrc_data_rsc_q)
    );
  DCT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_22_4194304_3_gen mdst_data_rsci (
      .we(mdst_data_rsc_we),
      .d(mdst_data_rsc_d),
      .wadr(mdst_data_rsc_wadr),
      .re(mdst_data_rsc_re),
      .q(mdst_data_rsc_q),
      .radr(mdst_data_rsc_radr),
      .radr_d(mdst_data_rsci_radr_d),
      .wadr_d(mdst_data_rsci_wadr_d),
      .d_d(mdst_data_rsci_d_d),
      .we_d(mdst_data_rsci_we_d),
      .re_d(mdst_data_rsci_re_d),
      .q_d(mdst_data_rsci_q_d)
    );
  DCT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_22_4194304_4_gen msrc_data_rsci (
      .we(msrc_data_rsc_we),
      .d(msrc_data_rsc_d),
      .wadr(msrc_data_rsc_wadr),
      .re(msrc_data_rsc_re),
      .q(msrc_data_rsc_q),
      .radr(msrc_data_rsc_radr),
      .radr_d(msrc_data_rsci_radr_d),
      .wadr_d(msrc_data_rsci_wadr_d),
      .d_d(msrc_data_rsci_d_d),
      .we_d(msrc_data_rsci_we_d),
      .re_d(msrc_data_rsci_re_d),
      .q_d(msrc_data_rsci_q_d)
    );
  DCT_core DCT_core_inst (
      .clk(clk),
      .rst(rst),
      .dst_rsc_dat(dst_rsc_dat),
      .dst_rsc_vld(dst_rsc_vld),
      .dst_rsc_rdy(dst_rsc_rdy),
      .src_rsc_dat(src_rsc_dat),
      .src_rsc_vld(src_rsc_vld),
      .src_rsc_rdy(src_rsc_rdy),
      .mdst_data_rsci_radr_d(mdst_data_rsci_radr_d),
      .mdst_data_rsci_wadr_d(mdst_data_rsci_wadr_d),
      .mdst_data_rsci_d_d(mdst_data_rsci_d_d),
      .mdst_data_rsci_we_d(mdst_data_rsci_we_d),
      .mdst_data_rsci_re_d(mdst_data_rsci_re_d),
      .mdst_data_rsci_q_d(mdst_data_rsci_q_d),
      .msrc_data_rsci_radr_d(msrc_data_rsci_radr_d),
      .msrc_data_rsci_wadr_d(msrc_data_rsci_wadr_d),
      .msrc_data_rsci_d_d(msrc_data_rsci_d_d),
      .msrc_data_rsci_we_d(msrc_data_rsci_we_d),
      .msrc_data_rsci_re_d(msrc_data_rsci_re_d),
      .msrc_data_rsci_q_d(msrc_data_rsci_q_d)
    );
endmodule



